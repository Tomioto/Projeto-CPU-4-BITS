CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
20
13 MT.Decode2bit
94 404 189 0 6 13
0 9 10 11 12 3 4
13 MT.Decode2bit
1 0 4224 0
0
2 U3
42 -9 56 -1
0
0
0
0
0
0
13

0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 1 0 0 0
1 U
5130 0 0
2
5.90094e-315 5.43451e-315
0
12 Hex Display~
7 729 80 0 16 19
10 2 31 32 33 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
2 Y1
-7 -38 7 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
391 0 0
2
5.90094e-315 5.43192e-315
0
14 Logic Display~
6 142 86 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 I7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
5.90094e-315 5.42933e-315
0
14 Logic Display~
6 162 86 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 I6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.90094e-315 5.42414e-315
0
14 Logic Display~
6 182 86 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 I5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.90094e-315 5.41896e-315
0
14 Logic Display~
6 202 86 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 I4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.90094e-315 5.41378e-315
0
14 Logic Display~
6 303 85 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.90094e-315 5.4086e-315
0
14 Logic Display~
6 283 85 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.90094e-315 5.40342e-315
0
14 Logic Display~
6 694 79 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.90094e-315 5.39824e-315
0
9 2-In AND~
219 472 299 0 3 22
0 12 8 17
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
972 0 0
2
5.90094e-315 5.39306e-315
0
9 2-In AND~
219 472 341 0 3 22
0 11 7 15
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
3472 0 0
2
5.90094e-315 5.38788e-315
0
9 2-In AND~
219 473 384 0 3 22
0 10 6 14
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9998 0 0
2
5.90094e-315 5.37752e-315
0
9 2-In AND~
219 473 426 0 3 22
0 9 5 16
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
3536 0 0
2
5.90094e-315 5.36716e-315
0
8 4-In OR~
219 602 357 0 5 22
0 17 15 14 16 2
0
0 0 96 0
4 4072
-14 -24 14 -16
3 U1A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 1 0
1 U
4597 0 0
2
5.90094e-315 5.3568e-315
0
8 Hex Key~
166 249 76 0 11 12
0 34 35 36 37 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD5
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
3835 0 0
2
5.90094e-315 5.34643e-315
0
8 Hex Key~
166 103 78 0 11 12
0 38 39 40 41 0 0 0 0 0
1 49
0
0 0 4640 0
0
2 I0
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
3670 0 0
2
5.90094e-315 5.32571e-315
0
8 Hex Key~
166 104 161 0 11 12
0 42 43 44 45 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I1
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
5616 0 0
2
5.90094e-315 5.30499e-315
0
8 Hex Key~
166 105 237 0 11 12
0 46 47 48 49 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I2
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9323 0 0
2
5.90094e-315 5.26354e-315
0
8 Hex Key~
166 104 311 0 11 12
0 50 51 52 53 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I3
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
317 0 0
2
5.90094e-315 0
0
9 MT.Mux4x1
94 484 532 0 1 15
0 0
9 MT.Mux4x1
2 0 4736 0
0
2 U4
50 0 64 8
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
3108 0 0
2
45193.9 0
0
44
5 0 2 0 0 8192 0 20 0 0 38 3
484 566
484 577
694 577
7 0 3 0 0 4352 0 20 0 0 40 2
432 541
283 541
6 0 4 0 0 4352 0 20 0 0 39 2
432 532
303 532
1 0 5 0 0 8192 0 20 0 0 44 3
448 507
448 502
142 502
2 0 6 0 0 8192 0 20 0 0 43 3
466 507
466 493
162 493
3 0 7 0 0 8192 0 20 0 0 42 3
502 507
502 485
182 485
4 0 8 0 0 8192 0 20 0 0 41 3
520 507
520 475
202 475
1 1 9 0 0 4224 0 1 13 0 0 3
359 213
359 417
449 417
2 1 10 0 0 4224 0 1 12 0 0 3
377 213
377 375
449 375
3 1 11 0 0 4224 0 1 11 0 0 3
413 213
413 332
448 332
4 1 12 0 0 4224 0 1 10 0 0 3
431 213
431 290
448 290
5 0 3 0 0 256 0 1 0 0 40 2
386 155
283 155
6 0 4 0 0 256 0 1 0 0 39 3
404 155
404 146
303 146
0 0 1 0 0 4256 0 0 0 0 0 2
724 215
908 215
0 0 1 0 0 32 0 0 0 0 0 2
766 179
766 285
0 0 1 0 0 32 0 0 0 0 0 2
839 179
839 285
0 0 1 0 0 32 0 0 0 0 0 6
729 179
908 179
908 285
724 285
724 179
729 179
0 0 1 0 0 32 0 0 0 0 0 2
744 36
685 36
0 0 1 0 0 32 0 0 0 0 0 2
233 41
312 41
0 0 1 0 0 32 0 0 0 0 0 2
89 41
210 41
0 0 13 0 0 8576 0 0 0 0 0 6
324 124
324 458
705 458
705 98
324 98
324 124
5 0 2 0 0 0 0 14 0 0 38 2
635 357
694 357
2 0 5 0 0 4096 0 13 0 0 44 2
449 435
142 435
2 0 6 0 0 0 0 12 0 0 43 2
449 393
162 393
2 0 7 0 0 0 0 11 0 0 42 2
448 350
182 350
2 0 8 0 0 0 0 10 0 0 41 2
448 308
202 308
3 3 14 0 0 12416 0 12 14 0 0 4
494 384
536 384
536 362
585 362
3 2 15 0 0 12416 0 11 14 0 0 4
493 341
536 341
536 353
585 353
3 4 16 0 0 8320 0 13 14 0 0 4
494 426
548 426
548 371
585 371
3 1 17 0 0 4224 0 10 14 0 0 4
493 299
548 299
548 344
585 344
0 0 3 0 0 256 0 0 0 0 40 3
251 105
251 140
283 140
0 0 4 0 0 256 0 0 0 0 39 3
257 105
257 124
303 124
0 0 5 0 0 0 0 0 0 0 44 3
114 340
114 347
142 347
0 0 6 0 0 0 0 0 0 0 43 3
114 267
114 276
162 276
0 0 7 0 0 0 0 0 0 0 42 3
113 190
113 201
182 201
0 0 8 0 0 0 0 0 0 0 41 3
112 107
112 120
202 120
1 0 2 0 0 0 0 2 0 0 38 3
738 104
738 131
694 131
1 0 2 0 0 4224 0 9 0 0 0 2
694 97
694 605
1 0 4 0 0 4480 0 7 0 0 0 2
303 103
303 604
1 0 3 0 0 4480 0 8 0 0 0 2
283 103
283 604
1 0 8 0 0 4224 0 6 0 0 0 2
202 104
202 604
1 0 7 0 0 4224 0 5 0 0 0 2
182 104
182 604
1 0 6 0 0 4224 0 4 0 0 0 2
162 104
162 605
1 0 5 0 0 4224 0 3 0 0 0 2
142 104
142 606
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
467 73 536 97
473 77 529 93
7 Mux.4x1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
127 19 172 43
133 23 165 39
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
689 13 742 37
695 17 735 33
5 Out's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
252 19 297 43
258 23 290 39
4 Ctrl
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
723 180 768 304
729 184 761 280
22 Dec.

 0
 1
 2
 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 96
770 180 911 304
776 184 904 280
96  Ctrl      Out's
S1  S0       Y
0   0       I0
0   1       I1
1   0       I2
1   1       I3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
