CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
15
12 Hex Display~
7 626 107 0 16 19
10 6 5 4 3 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3751 0 0
2
45194.8 13
0
14 Logic Display~
6 133 111 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4292 0 0
2
45194.8 12
0
14 Logic Display~
6 153 111 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6118 0 0
2
45194.8 11
0
14 Logic Display~
6 591 112 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
45194.8 10
0
14 Logic Display~
6 531 112 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
45194.8 9
0
14 Logic Display~
6 551 112 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
45194.8 8
0
14 Logic Display~
6 571 112 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 M1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3976 0 0
2
45194.8 7
0
9 Inverter~
13 177 168 0 2 22
0 8 10
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U2B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
7634 0 0
2
45194.8 6
0
9 Inverter~
13 201 169 0 2 22
0 7 9
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U2A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
523 0 0
2
45194.8 5
0
9 2-In AND~
219 255 218 0 3 22
0 10 9 6
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
6748 0 0
2
45194.8 4
0
9 2-In AND~
219 254 253 0 3 22
0 10 7 5
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
6901 0 0
2
45194.8 3
0
9 2-In AND~
219 254 288 0 3 22
0 8 9 4
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
842 0 0
2
45194.8 2
0
9 2-In AND~
219 254 324 0 3 22
0 8 7 3
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3277 0 0
2
45194.8 1
0
8 Hex Key~
166 101 102 0 11 12
0 7 8 11 12 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
4212 0 0
2
45194.8 0
0
13 MT.Decode2bit
94 365 423 0 1 13
0 0
13 MT.Decode2bit
1 0 4736 0
0
2 U3
42 -9 56 -1
0
0
0
0
0
0
13

0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 0 0 0 0
1 U
4720 0 0
2
45193.9 0
0
41
0 0 -1 0 0 272 0 0 0 0 0 5
120 128
608 128
608 374
120 374
120 128
1 0 -1 0 0 16 0 15 0 0 19 5
320 447
320 466
526 466
526 433
531 433
2 0 -1 0 0 16 0 15 0 0 18 5
338 447
338 461
546 461
546 429
551 429
3 0 -1 0 0 16 0 15 0 0 17 5
374 447
374 456
566 456
566 440
571 440
4 0 -1 0 0 16 0 15 0 0 16 3
392 447
392 451
591 451
5 0 -1 0 0 16 0 15 0 0 23 2
347 389
133 389
6 0 -1 0 0 16 0 15 0 0 22 3
365 389
365 381
153 381
1 0 -1 0 0 16 0 13 0 0 23 2
230 315
133 315
2 0 -1 0 0 16 0 13 0 0 22 2
230 333
153 333
1 0 -1 0 0 16 0 12 0 0 23 2
230 279
133 279
2 0 -1 0 0 16 0 11 0 0 22 2
230 262
153 262
1 0 -1 0 0 16 0 1 0 0 16 3
635 131
635 170
591 170
2 0 -1 0 0 16 0 1 0 0 17 3
629 131
629 158
571 158
3 0 -1 0 0 16 0 1 0 0 18 3
623 131
623 147
551 147
4 0 -1 0 0 16 0 1 0 0 19 3
617 131
617 139
531 139
1 0 -1 0 0 16 0 4 0 0 0 2
591 130
591 471
1 0 -1 0 0 16 0 7 0 0 0 2
571 130
571 472
1 0 -1 0 0 16 0 6 0 0 0 2
551 130
551 472
1 0 -1 0 0 16 0 5 0 0 0 2
531 130
531 472
1 0 -1 0 0 16 0 8 0 0 23 3
180 150
180 141
133 141
1 0 -1 0 0 16 0 9 0 0 22 3
204 151
204 133
153 133
1 0 -1 0 0 16 0 3 0 0 0 2
153 129
153 473
1 0 -1 0 0 16 0 2 0 0 0 2
133 129
133 473
0 0 -1 0 0 48 0 0 0 0 0 2
641 63
521 63
0 0 -1 0 0 48 0 0 0 0 0 2
83 62
161 62
0 0 -1 0 0 48 0 0 0 0 0 2
628 233
841 233
0 0 -1 0 0 48 0 0 0 0 0 2
668 213
668 303
0 0 -1 0 0 48 0 0 0 0 0 2
727 213
727 303
0 0 -1 0 0 48 0 0 0 0 0 5
628 213
841 213
841 303
628 303
628 213
3 0 -1 0 0 16 0 13 0 0 0 2
275 324
531 324
3 0 -1 0 0 16 0 12 0 0 0 2
275 288
551 288
3 0 -1 0 0 16 0 11 0 0 0 2
275 253
571 253
3 0 -1 0 0 16 0 10 0 0 0 2
276 218
591 218
2 0 -1 0 0 272 0 12 0 0 39 2
230 297
204 297
1 0 -1 0 0 272 0 11 0 0 38 2
230 244
180 244
2 0 -1 0 0 272 0 10 0 0 39 2
231 227
204 227
1 0 -1 0 0 272 0 10 0 0 38 2
231 209
180 209
2 0 -1 0 0 272 0 8 0 0 0 2
180 186
180 368
2 0 -1 0 0 272 0 9 0 0 0 2
204 187
204 368
0 0 -1 0 0 16 0 0 0 0 0 3
103 130
103 179
133 179
0 0 -1 0 0 16 0 0 0 0 0 3
109 130
109 167
153 167
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
627 212 672 316
633 216 665 296
16 Dec.
0
1
2
3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 105
668 214 841 318
674 218 834 298
105 S1 S0    M3 M2 M1 M0
0  0     0  0  0  1
0  1     0  0  1  0 
1  0     0  1  0  0
1  1     1  0  0  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
308 103 401 127
314 107 394 123
10 Decode2bit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
99 39 144 63
105 43 137 59
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
555 40 608 64
561 44 601 60
5 Out's
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
