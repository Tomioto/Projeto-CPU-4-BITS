CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
8912914 0
0
6 Title:
5 Name:
0
0
0
19
10 2-In NAND~
219 725 412 0 1 22
0 0
0
0 0 96 270
6 74LS00
-14 -24 28 -16
3 U1D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3108 0 0
2
45193.1 0
0
10 2-In NAND~
219 684 412 0 1 22
0 0
0
0 0 96 270
6 74LS00
-14 -24 28 -16
3 U1C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
4299 0 0
2
45193.1 0
0
10 2-In NAND~
219 643 412 0 1 22
0 0
0
0 0 96 270
6 74LS00
-14 -24 28 -16
3 U1B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
9672 0 0
2
45193.1 0
0
10 2-In NAND~
219 600 413 0 1 22
0 0
0
0 0 96 270
6 74LS00
-14 -24 28 -16
3 U1A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
7876 0 0
2
45193.1 0
0
14 Logic Display~
6 924 447 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
45193.1 0
0
14 Logic Display~
6 944 447 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
45193.1 1
0
14 Logic Display~
6 965 447 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
45193.1 2
0
14 Logic Display~
6 986 447 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
45193.1 3
0
8 Hex Key~
166 328 101 0 11 12
0 13 14 15 16 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7678 0 0
2
45193.1 4
0
14 Logic Display~
6 449 87 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
45193.1 5
0
14 Logic Display~
6 428 87 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
45193.1 6
0
14 Logic Display~
6 407 87 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
45193.1 7
0
14 Logic Display~
6 387 87 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
45193.1 8
0
14 Logic Display~
6 267 89 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
45193.1 9
0
14 Logic Display~
6 246 89 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
45193.1 10
0
14 Logic Display~
6 223 89 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
45193.1 11
0
14 Logic Display~
6 201 89 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
45193.1 12
0
8 Hex Key~
166 160 104 0 11 12
0 13 14 15 16 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9424 0 0
2
45193.1 13
0
12 Hex Display~
7 1044 462 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusY
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9968 0 0
2
45193.1 14
0
58
0 0 0 0 0 0 0 0 0 0 0 2
691 91
780 91
3 0 0 0 0 0 0 1 0 0 34 2
726 438
726 510
3 0 0 0 0 0 0 2 0 0 32 2
685 438
685 522
3 0 0 0 0 0 0 3 0 0 33 2
644 438
644 535
3 0 0 0 0 0 0 4 0 0 31 2
601 439
601 548
0 0 8 0 0 272 0 0 0 0 0 6
27 272
27 336
83 336
83 266
27 266
27 272
0 0 8 0 0 256 0 0 0 0 0 6
27 168
27 232
83 232
83 162
27 162
27 168
0 0 0 0 0 32 0 0 0 0 0 2
625 58
625 119
0 0 0 0 0 32 0 0 0 0 0 2
523 81
795 81
0 0 0 0 0 32 0 0 0 0 0 5
523 58
795 58
795 119
523 119
523 58
0 0 0 0 0 256 0 0 0 0 0 5
501 157
501 568
778 568
778 153
501 153
1 0 0 0 0 0 0 1 0 0 58 2
735 387
735 282
2 0 0 0 0 0 0 1 0 0 54 2
717 387
717 176
1 0 0 0 0 0 0 2 0 0 57 4
694 387
694 311
671 311
671 296
2 0 0 0 0 0 0 2 0 0 53 4
676 387
676 205
653 205
653 190
1 0 0 0 0 0 0 3 0 0 56 4
653 387
653 325
608 325
608 310
2 0 0 0 0 0 0 3 0 0 52 4
635 387
635 219
590 219
590 204
1 0 0 0 0 0 0 4 0 0 55 4
610 388
610 338
541 338
541 323
2 0 0 0 0 0 0 4 0 0 51 4
592 388
592 232
523 232
523 217
0 0 1 0 0 32 0 0 0 0 0 2
913 416
1062 416
0 0 1 0 0 4256 0 0 0 0 0 2
143 60
459 60
1 0 2 0 0 4096 0 19 0 0 34 2
1053 486
1053 510
2 0 3 0 0 4096 0 19 0 0 32 2
1047 486
1047 522
3 0 4 0 0 4096 0 19 0 0 33 2
1041 486
1041 535
4 0 5 0 0 4096 0 19 0 0 31 2
1035 486
1035 548
1 0 2 0 0 4096 0 8 0 0 34 2
986 465
986 510
1 0 3 0 0 4096 0 7 0 0 32 2
965 465
965 522
1 0 4 0 0 4096 0 6 0 0 33 2
944 465
944 535
1 0 5 0 0 4096 0 5 0 0 31 2
924 465
924 548
0 0 6 0 0 12672 0 0 0 0 0 6
1081 499
1081 563
1138 563
1138 490
1081 490
1081 499
0 0 5 0 0 4224 0 0 0 0 0 2
56 548
1112 548
0 0 3 0 0 4224 0 0 0 0 0 2
57 522
1113 522
0 0 4 0 0 4224 0 0 0 0 0 2
58 535
1112 535
0 0 2 0 0 4224 0 0 0 0 0 2
57 510
1113 510
1 0 9 0 0 4096 0 10 0 0 58 2
449 105
449 282
1 0 10 0 0 4096 0 11 0 0 57 2
428 105
428 296
1 0 11 0 0 4096 0 12 0 0 56 2
407 105
407 310
1 0 12 0 0 4096 0 13 0 0 55 2
387 105
387 323
1 0 13 0 0 4096 0 9 0 0 54 2
337 125
337 176
2 0 14 0 0 4096 0 9 0 0 53 2
331 125
331 190
3 0 15 0 0 4096 0 9 0 0 52 2
325 125
325 204
4 0 16 0 0 4096 0 9 0 0 51 2
319 125
319 217
1 0 13 0 0 4096 0 14 0 0 54 2
267 107
267 176
1 0 14 0 0 4096 0 15 0 0 53 2
246 107
246 190
1 0 15 0 0 4096 0 16 0 0 52 2
223 107
223 204
1 0 16 0 0 4096 0 17 0 0 51 2
201 107
201 217
1 0 13 0 0 0 0 18 0 0 54 2
169 128
169 176
2 0 14 0 0 0 0 18 0 0 53 2
163 128
163 190
3 0 15 0 0 0 0 18 0 0 52 2
157 128
157 204
4 0 16 0 0 0 0 18 0 0 51 2
151 128
151 217
0 0 16 0 0 4224 0 0 0 0 0 2
54 217
937 217
0 0 15 0 0 4224 0 0 0 0 0 2
55 204
937 204
0 0 14 0 0 4224 0 0 0 0 0 2
55 190
938 190
0 0 13 0 0 4224 0 0 0 0 0 2
53 176
939 176
0 0 12 0 0 4224 0 0 0 0 0 2
55 323
938 323
0 0 11 0 0 4224 0 0 0 0 0 2
56 310
938 310
0 0 10 0 0 4224 0 0 0 0 0 2
56 296
939 296
0 0 9 0 0 4224 0 0 0 0 0 2
54 282
940 282
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
592 35 685 59
598 39 678 55
10 Nand.4bits
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
591 129 684 153
597 133 677 149
10 Nand.4bits
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 60
521 59 790 123
527 63 783 111
60    In's            Out's

 BusA, BusB   BusY = BusA . BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1080 467 1125 491
1086 471 1118 487
4 BusY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
32 138 77 162
38 142 70 158
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
34 244 79 268
40 248 72 264
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
266 36 311 60
272 40 304 56
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
960 392 1013 416
966 396 1006 412
5 Out's
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
