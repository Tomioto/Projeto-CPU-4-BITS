CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 75 1364 626
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 171 457 268
8912914 0
0
6 Title:
5 Name:
0
0
0
21
14 Logic Display~
6 250 424 0 1 2
10 0
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 Ts3
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5130 0 0
2
45193.9 0
0
7 Ground~
168 791 437 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
391 0 0
2
45193.9 0
0
14 Logic Display~
6 924 447 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Z3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
45193.9 0
0
14 Logic Display~
6 944 447 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Z2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
45193.9 1
0
14 Logic Display~
6 965 447 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Z1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
45193.9 2
0
14 Logic Display~
6 986 447 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Z0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
45193.9 3
0
8 Hex Key~
166 328 101 0 11 12
0 13 14 15 16 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8901 0 0
2
45193.9 4
0
14 Logic Display~
6 449 87 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
45193.9 5
0
14 Logic Display~
6 428 87 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
45193.9 6
0
14 Logic Display~
6 407 87 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
45193.9 7
0
14 Logic Display~
6 387 87 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
45193.9 8
0
14 Logic Display~
6 267 89 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
45193.9 9
0
14 Logic Display~
6 246 89 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
45193.9 10
0
14 Logic Display~
6 223 89 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
45193.9 11
0
14 Logic Display~
6 201 89 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
45193.9 12
0
8 Hex Key~
166 160 104 0 11 12
0 13 14 15 16 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3670 0 0
2
45193.9 13
0
12 Hex Display~
7 1044 462 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5616 0 0
2
45193.9 14
0
10 MT.Sub1bit
94 335 426 0 1 11
0 0
10 MT.Sub1bit
1 0 4736 0
0
2 U1
56 -32 70 -24
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
9323 0 0
2
45193.9 0
0
10 MT.Sub1bit
94 461 425 0 1 11
0 0
10 MT.Sub1bit
2 0 4736 0
0
2 U2
56 -32 70 -24
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
317 0 0
2
45193.9 0
0
10 MT.Sub1bit
94 586 424 0 1 11
0 0
10 MT.Sub1bit
3 0 4736 0
0
2 U3
56 -32 70 -24
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
3108 0 0
2
45193.9 0
0
10 MT.Sub1bit
94 711 423 0 1 11
0 0
10 MT.Sub1bit
4 0 4736 0
0
2 U4
56 -32 70 -24
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
4299 0 0
2
45193.9 0
0
61
1 2 0 0 0 0 0 1 18 0 0 2
265 427
279 427
1 0 0 0 0 0 0 21 0 0 35 2
711 453
711 510
1 0 0 0 0 0 0 20 0 0 33 2
586 454
586 522
1 0 0 0 0 0 0 19 0 0 34 2
461 455
461 535
1 0 0 0 0 0 0 18 0 0 32 2
335 456
335 548
5 0 0 0 0 0 0 21 0 0 61 2
734 394
734 282
4 0 0 0 0 0 0 21 0 0 57 2
689 395
689 176
5 0 0 0 0 0 0 20 0 0 60 2
609 395
609 296
4 0 0 0 0 0 0 20 0 0 56 2
564 396
564 190
5 0 0 0 0 0 0 19 0 0 59 2
484 396
484 310
4 0 0 0 0 0 0 19 0 0 55 2
439 397
439 204
5 0 0 0 0 0 0 18 0 0 58 2
358 397
358 323
4 0 0 0 0 0 0 18 0 0 54 2
313 398
313 217
3 1 0 0 0 0 0 21 2 0 0 3
768 423
791 423
791 431
3 2 0 0 0 0 0 20 21 0 0 2
643 424
655 424
3 2 0 0 0 0 0 19 20 0 0 2
518 425
530 425
3 2 0 0 0 0 0 18 19 0 0 2
392 426
405 426
0 0 1 0 0 4128 0 0 0 0 0 2
541 73
798 73
0 0 1 0 0 32 0 0 0 0 0 2
635 59
635 96
0 0 1 0 0 4128 0 0 0 0 0 5
538 59
798 59
798 96
538 96
538 59
0 0 1 0 0 32 0 0 0 0 0 2
913 416
1062 416
0 0 1 0 0 4256 0 0 0 0 0 2
143 60
459 60
1 0 2 0 0 4096 0 17 0 0 35 2
1053 486
1053 510
2 0 3 0 0 4096 0 17 0 0 33 2
1047 486
1047 522
3 0 4 0 0 4096 0 17 0 0 34 2
1041 486
1041 535
4 0 5 0 0 4096 0 17 0 0 32 2
1035 486
1035 548
1 0 2 0 0 4096 0 6 0 0 35 2
986 465
986 510
1 0 3 0 0 4096 0 5 0 0 33 2
965 465
965 522
1 0 4 0 0 4096 0 4 0 0 34 2
944 465
944 535
1 0 5 0 0 4096 0 3 0 0 32 2
924 465
924 548
0 0 6 0 0 12672 0 0 0 0 0 6
1081 499
1081 563
1138 563
1138 490
1081 490
1081 499
0 0 5 0 0 4224 0 0 0 0 0 2
56 548
1112 548
0 0 3 0 0 4224 0 0 0 0 0 2
57 522
1113 522
0 0 4 0 0 4224 0 0 0 0 0 2
58 535
1112 535
0 0 2 0 0 4224 0 0 0 0 0 2
57 510
1113 510
0 0 7 0 0 12672 0 0 0 0 0 6
918 273
918 337
975 337
975 264
918 264
918 273
0 0 8 0 0 12672 0 0 0 0 0 6
917 164
917 230
975 230
975 158
917 158
917 164
1 0 9 0 0 4096 0 8 0 0 61 2
449 105
449 282
1 0 10 0 0 4096 0 9 0 0 60 2
428 105
428 296
1 0 11 0 0 4096 0 10 0 0 59 2
407 105
407 310
1 0 12 0 0 4096 0 11 0 0 58 2
387 105
387 323
1 0 13 0 0 4096 0 7 0 0 57 2
337 125
337 176
2 0 14 0 0 4096 0 7 0 0 56 2
331 125
331 190
3 0 15 0 0 4096 0 7 0 0 55 2
325 125
325 204
4 0 16 0 0 4096 0 7 0 0 54 2
319 125
319 217
1 0 13 0 0 4096 0 12 0 0 57 2
267 107
267 176
1 0 14 0 0 4096 0 13 0 0 56 2
246 107
246 190
1 0 15 0 0 4096 0 14 0 0 55 2
223 107
223 204
1 0 16 0 0 4096 0 15 0 0 54 2
201 107
201 217
1 0 13 0 0 0 0 16 0 0 57 2
169 128
169 176
2 0 14 0 0 0 0 16 0 0 56 2
163 128
163 190
3 0 15 0 0 0 0 16 0 0 55 2
157 128
157 204
4 0 16 0 0 0 0 16 0 0 54 2
151 128
151 217
0 0 16 0 0 4224 0 0 0 0 0 2
54 217
937 217
0 0 15 0 0 4224 0 0 0 0 0 2
55 204
937 204
0 0 14 0 0 4224 0 0 0 0 0 2
55 190
938 190
0 0 13 0 0 4224 0 0 0 0 0 2
53 176
939 176
0 0 12 0 0 4224 0 0 0 0 0 2
55 323
938 323
0 0 11 0 0 4224 0 0 0 0 0 2
56 310
938 310
0 0 10 0 0 4224 0 0 0 0 0 2
56 296
939 296
0 0 9 0 0 4224 0 0 0 0 0 2
54 282
940 282
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
916 135 961 159
922 139 954 155
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
266 36 311 60
272 40 304 56
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
960 392 1013 416
966 396 1006 412
5 Out's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1080 467 1125 491
1086 471 1118 487
4 BusZ
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
917 242 962 266
923 246 955 262
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 58
531 55 800 99
537 59 793 91
58    In's            Out's
 BusA, BusB   Busz = BusA + BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
539 122 728 146
545 126 721 142
22 * Subtrator Aritm�tico
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
606 34 691 58
612 38 684 54
9 Sub.4bits
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
