CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
8912914 0
0
6 Title:
5 Name:
0
0
0
12
9 2-In AND~
219 236 365 0 3 22
0 4 5 8
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 5 0
1 U
631 0 0
2
45189.8 0
0
8 2-In OR~
219 412 361 0 3 22
0 7 8 2
0
0 0 624 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
9466 0 0
2
45189.8 0
0
9 2-In AND~
219 319 286 0 3 22
0 9 6 7
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 5 0
1 U
3266 0 0
2
45189.8 0
0
9 2-In XOR~
219 223 220 0 3 22
0 4 5 9
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7693 0 0
2
45189.8 0
0
9 2-In XOR~
219 309 160 0 3 22
0 6 9 3
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3723 0 0
2
45189.8 0
0
14 Logic Display~
6 501 78 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Ts
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3440 0 0
2
45189.8 0
0
14 Logic Display~
6 526 78 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 W
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6263 0 0
2
45189.8 0
0
14 Logic Display~
6 185 83 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Te
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4900 0 0
2
45189.8 0
0
14 Logic Display~
6 162 83 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8783 0 0
2
45189.8 0
0
14 Logic Display~
6 139 83 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3221 0 0
2
45189.8 0
0
12 Hex Display~
7 581 91 0 18 19
10 3 2 11 12 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
3215 0 0
2
45189.8 0
0
8 Hex Key~
166 81 96 0 11 12
0 6 5 4 13 0 0 0 0 0
4 52
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
7903 0 0
2
45189.8 0
0
30
0 0 1 0 0 4128 0 0 0 0 0 2
626 183
870 183
0 0 1 0 0 32 0 0 0 0 0 5
622 360
832 360
832 401
622 401
622 360
0 0 1 0 0 32 0 0 0 0 0 2
820 159
820 318
0 0 1 0 0 32 0 0 0 0 0 2
750 159
750 318
0 0 1 0 0 32 0 0 0 0 0 2
671 159
671 318
0 0 1 0 0 32 0 0 0 0 0 5
626 159
870 159
870 318
626 318
626 159
0 0 1 0 0 4256 0 0 0 0 0 2
129 255
538 255
2 0 2 0 0 8192 0 11 0 0 27 3
584 115
584 133
501 133
1 0 3 0 0 8192 0 11 0 0 26 3
590 115
590 143
526 143
3 0 4 0 0 8192 0 12 0 0 30 3
78 120
78 141
139 141
2 0 5 0 0 8192 0 12 0 0 29 3
84 120
84 129
162 129
1 0 6 0 0 4096 0 12 0 0 28 2
90 120
185 120
3 0 2 0 0 0 0 2 0 0 27 2
445 361
501 361
3 0 3 0 0 4096 0 5 0 0 26 2
342 160
526 160
3 1 7 0 0 8320 0 3 2 0 0 4
340 286
392 286
392 352
399 352
3 2 8 0 0 4224 0 1 2 0 0 4
257 365
390 365
390 370
399 370
2 0 5 0 0 0 0 1 0 0 29 2
212 374
162 374
1 0 4 0 0 4096 0 1 0 0 30 2
212 356
139 356
2 0 6 0 0 4096 0 3 0 0 28 2
295 295
185 295
2 0 5 0 0 0 0 4 0 0 29 2
207 229
162 229
1 0 4 0 0 0 0 4 0 0 30 2
207 211
139 211
0 1 9 0 0 4480 0 0 3 23 0 3
282 220
282 277
295 277
3 2 9 0 0 0 0 4 5 0 0 4
256 220
283 220
283 169
293 169
1 0 6 0 0 0 0 5 0 0 28 2
293 151
185 151
0 0 10 0 0 12672 0 0 0 0 0 5
123 99
548 99
548 456
118 456
118 99
1 0 3 0 0 4224 0 7 0 0 0 2
526 96
526 437
1 0 2 0 0 4224 0 6 0 0 0 2
501 96
501 438
1 0 6 0 0 4224 0 8 0 0 0 2
185 101
185 438
1 0 5 0 0 4224 0 9 0 0 0 2
162 101
162 439
1 0 4 0 0 4224 0 10 0 0 0 2
139 101
139 440
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 45
622 361 835 405
628 365 828 397
45 W = A (+) B (+) Te
Ts = A.B + Te . (A (+) B)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
835 183 856 347
841 187 849 315
22 0
1
2
3
4
5
6
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
637 181 658 345
643 185 651 313
22 0
1
2
3
4
5
6
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
825 163 870 187
831 167 863 183
4 Dec.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
625 163 670 187
631 166 663 182
4 Dec.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 52
765 165 810 349
771 169 803 313
52 Ts W
0  0
0  1
0  1
1  0
0  1
1  0
1  0
1  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 63
677 163 738 347
683 167 731 311
63 A B Te
0 0 0 
0 0 1
0 1 0
0 1 1
1 0 0
1 0 1
1 1 0
1 1 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
