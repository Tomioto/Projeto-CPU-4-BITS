CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
22
10 MT.Add1bit
94 763 419 0 1 11
0 0
10 MT.Add1bit
9 0 4224 0
0
2 U4
68 -36 82 -28
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
4597 0 0
2
45194.8 56
0
10 MT.Add1bit
94 621 420 0 1 11
0 0
10 MT.Add1bit
8 0 4224 0
0
2 U3
68 -36 82 -28
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
3835 0 0
2
45194.8 43
0
10 MT.Add1bit
94 478 421 0 1 11
0 0
10 MT.Add1bit
7 0 4224 0
0
2 U2
68 -36 82 -28
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
3670 0 0
2
45194.8 30
0
10 MT.Add1bit
94 335 422 0 1 11
0 0
10 MT.Add1bit
6 0 4224 0
0
2 U1
68 -36 82 -28
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
5616 0 0
2
45194.8 17
0
12 Hex Display~
7 1017 452 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9323 0 0
2
45194.8 16
0
14 Logic Display~
6 174 79 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
45194.8 15
0
14 Logic Display~
6 196 79 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
45194.8 14
0
14 Logic Display~
6 219 79 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
45194.8 13
0
14 Logic Display~
6 240 79 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9672 0 0
2
45194.8 12
0
14 Logic Display~
6 360 77 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
45194.8 11
0
14 Logic Display~
6 380 77 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
45194.8 10
0
14 Logic Display~
6 401 77 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
45194.8 9
0
14 Logic Display~
6 422 77 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
45194.8 8
0
14 Logic Display~
6 959 437 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 W0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
45194.8 7
0
14 Logic Display~
6 938 437 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 W1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
45194.8 6
0
14 Logic Display~
6 917 437 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 W2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
45194.8 5
0
14 Logic Display~
6 897 437 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 W3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3178 0 0
2
45194.8 4
0
7 Ground~
168 852 432 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3409 0 0
2
45194.8 3
0
14 Logic Display~
6 254 403 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 Ts3
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3951 0 0
2
45194.8 2
0
8 Hex Key~
166 133 87 0 11 12
0 13 14 15 16 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8885 0 0
2
45194.8 1
0
8 Hex Key~
166 301 87 0 11 12
0 13 14 15 16 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
3780 0 0
2
45194.8 0
0
10 MT.Add4bit
94 103 413 0 1 25
0 0
10 MT.Add4bit
1 0 4736 0
0
2 U5
42 0 56 8
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
9265 0 0
2
45193.9 0
0
73
1 0 -1 0 0 0 0 1 0 0 47 2
763 444
763 500
1 0 -1 0 0 0 0 2 0 0 45 2
621 445
621 512
1 0 -1 0 0 0 0 3 0 0 46 2
478 446
478 525
1 0 -1 0 0 0 0 4 0 0 44 2
335 447
335 538
5 0 -1 0 0 0 0 1 0 0 73 2
798 386
798 272
4 0 -1 0 0 0 0 1 0 0 69 2
735 386
735 166
5 0 -1 0 0 0 0 2 0 0 72 2
656 387
656 286
4 0 -1 0 0 0 0 2 0 0 68 2
593 387
593 180
5 0 -1 0 0 0 0 3 0 0 71 2
513 388
513 300
4 0 -1 0 0 0 0 3 0 0 67 2
450 388
450 194
5 0 -1 0 0 0 0 4 0 0 70 2
370 389
370 313
4 0 -1 0 0 0 0 4 0 0 66 2
307 389
307 207
4 0 -1 0 0 0 0 22 0 0 47 2
130 446
130 500
3 0 -1 0 0 0 0 22 0 0 45 2
112 446
112 512
2 0 -1 0 0 0 0 22 0 0 46 2
76 446
76 525
1 0 -1 0 0 0 0 22 0 0 44 2
58 446
58 538
9 0 -1 0 0 0 0 22 0 0 70 2
103 389
103 313
10 0 -1 0 0 0 0 22 0 0 71 2
112 389
112 300
11 0 -1 0 0 0 0 22 0 0 72 4
121 389
121 291
122 291
122 286
12 0 -1 0 0 0 0 22 0 0 73 2
131 389
131 272
5 0 -1 0 0 0 0 22 0 0 66 2
58 389
58 207
6 0 -1 0 0 0 0 22 0 0 67 2
67 389
67 194
7 0 -1 0 0 0 0 22 0 0 68 2
77 389
77 180
8 0 -1 0 0 0 0 22 0 0 69 2
86 389
86 166
1 2 -1 0 0 0 0 19 4 0 0 3
254 421
254 423
271 423
3 1 -1 0 0 0 0 1 18 0 0 3
833 419
852 419
852 426
3 2 -1 0 0 0 0 2 1 0 0 2
691 420
699 420
3 2 -1 0 0 0 0 3 2 0 0 2
548 421
557 421
3 2 -1 0 0 0 0 4 3 0 0 2
405 422
414 422
0 0 -1 0 0 32 0 0 0 0 0 2
514 63
771 63
0 0 -1 0 0 32 0 0 0 0 0 2
608 49
608 86
0 0 -1 0 0 32 0 0 0 0 0 5
511 49
771 49
771 86
511 86
511 49
0 0 -1 0 0 32 0 0 0 0 0 2
886 406
1035 406
0 0 -1 0 0 32 0 0 0 0 0 2
116 50
432 50
1 0 -1 0 0 0 0 5 0 0 47 2
1026 476
1026 500
2 0 -1 0 0 0 0 5 0 0 45 2
1020 476
1020 512
3 0 -1 0 0 0 0 5 0 0 46 2
1014 476
1014 525
4 0 -1 0 0 0 0 5 0 0 44 2
1008 476
1008 538
1 0 -1 0 0 0 0 14 0 0 47 2
959 455
959 500
1 0 -1 0 0 0 0 15 0 0 45 2
938 455
938 512
1 0 -1 0 0 0 0 16 0 0 46 2
917 455
917 525
1 0 -1 0 0 0 0 17 0 0 44 2
897 455
897 538
0 0 -1 0 0 256 0 0 0 0 0 6
1054 489
1054 553
1111 553
1111 480
1054 480
1054 489
0 0 -1 0 0 0 0 0 0 0 0 2
29 538
1085 538
0 0 -1 0 0 0 0 0 0 0 0 2
30 512
1086 512
0 0 -1 0 0 0 0 0 0 0 0 2
31 525
1085 525
0 0 -1 0 0 0 0 0 0 0 0 2
30 500
1086 500
0 0 -1 0 0 256 0 0 0 0 0 6
891 263
891 327
948 327
948 254
891 254
891 263
0 0 -1 0 0 256 0 0 0 0 0 6
890 154
890 220
948 220
948 148
890 148
890 154
1 0 -1 0 0 0 0 13 0 0 73 2
422 95
422 272
1 0 -1 0 0 0 0 12 0 0 72 2
401 95
401 286
1 0 -1 0 0 0 0 11 0 0 71 2
380 95
380 300
1 0 -1 0 0 0 0 10 0 0 70 2
360 95
360 313
0 0 -1 0 0 0 0 0 0 0 69 2
310 115
310 166
0 0 -1 0 0 0 0 0 0 0 68 2
304 115
304 180
0 0 -1 0 0 0 0 0 0 0 67 2
298 115
298 194
0 0 -1 0 0 0 0 0 0 0 66 2
292 115
292 207
1 0 -1 0 0 0 0 9 0 0 69 2
240 97
240 166
1 0 -1 0 0 0 0 8 0 0 68 2
219 97
219 180
1 0 -1 0 0 0 0 7 0 0 67 2
196 97
196 194
1 0 -1 0 0 0 0 6 0 0 66 2
174 97
174 207
0 0 -1 0 0 0 0 0 0 0 69 3
141 115
142 115
142 166
0 0 -1 0 0 0 0 0 0 0 68 3
135 115
136 115
136 180
0 0 -1 0 0 0 0 0 0 0 67 3
129 115
130 115
130 194
0 0 -1 0 0 0 0 0 0 0 66 3
123 115
124 115
124 207
0 0 -1 0 0 0 0 0 0 0 0 2
27 207
910 207
0 0 -1 0 0 0 0 0 0 0 0 2
28 194
910 194
0 0 -1 0 0 0 0 0 0 0 0 2
28 180
911 180
0 0 -1 0 0 0 0 0 0 0 0 2
26 166
912 166
0 0 -1 0 0 0 0 0 0 0 0 2
26 313
911 313
0 0 -1 0 0 0 0 0 0 0 0 2
29 300
911 300
0 0 -1 0 0 0 0 0 0 0 0 2
29 286
912 286
0 0 -1 0 0 0 0 0 0 0 0 2
26 272
913 272
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1053 457 1098 481
1059 461 1091 477
4 BusW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
889 125 934 149
895 129 927 145
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
890 232 935 256
896 236 928 252
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
239 26 284 50
245 30 277 46
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
933 382 986 406
939 386 979 402
5 Out's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
512 112 661 156
518 116 654 148
17 * Soma Aritm�tica
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 58
504 45 773 89
510 49 766 81
58    In's            Out's
 BusA, BusB   BusW = BusA + BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
579 24 656 48
585 28 649 44
8 Add4bits
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
