CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 75 1364 626
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 171 457 268
8912914 0
0
6 Title:
5 Name:
0
0
0
19
8 4-In OR~
219 586 365 0 5 22
0 11 9 8 10 3
0
0 0 96 0
4 4072
-14 -24 14 -16
3 U3A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
9672 0 0
2
5.90094e-315 0
0
9 2-In AND~
219 461 434 0 3 22
0 14 4 10
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 4 2 0
1 U
7876 0 0
2
5.90094e-315 0
0
9 2-In AND~
219 461 392 0 3 22
0 15 5 8
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 3 2 0
1 U
6369 0 0
2
5.90094e-315 0
0
9 2-In AND~
219 460 349 0 3 22
0 16 6 9
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 2 2 0
1 U
9172 0 0
2
5.90094e-315 0
0
9 2-In AND~
219 460 307 0 3 22
0 17 7 11
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 512 4 1 2 0
1 U
7100 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 682 87 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 Y
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 271 93 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.90094e-315 5.26354e-315
0
14 Logic Display~
6 291 93 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.90094e-315 0
0
8 Hex Key~
166 236 89 0 11 12
0 13 12 18 19 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD5
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
3178 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 190 94 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 I0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3409 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 170 94 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 I1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 150 94 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 I2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8885 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 130 94 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 I3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3780 0 0
2
5.90094e-315 0
0
8 Hex Key~
166 93 324 0 11 12
0 4 20 21 22 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I3
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9265 0 0
2
5.90094e-315 0
0
8 Hex Key~
166 93 251 0 11 12
0 5 23 24 25 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I2
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9442 0 0
2
5.90094e-315 0
0
8 Hex Key~
166 92 174 0 11 12
0 6 26 27 28 0 0 0 0 0
0 48
0
0 0 4640 0
0
2 I1
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9424 0 0
2
5.90094e-315 0
0
8 Hex Key~
166 91 91 0 11 12
0 7 29 30 31 0 0 0 0 0
1 49
0
0 0 4640 0
0
2 I0
-7 -34 7 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9968 0 0
2
5.90094e-315 0
0
12 Hex Display~
7 717 88 0 16 19
10 3 32 33 34 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
1 Y
-4 -38 3 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
9281 0 0
2
5.90094e-315 0
0
13 MT.Decode2bit
94 392 197 0 1 13
0 0
13 MT.Decode2bit
1 0 4224 0
0
2 U1
42 -9 56 -1
0
0
0
0
0
0
13

0 0 0 0 0 0 0 0 0 0
0 0 0 0
0 0 0 0 0 0 0 0
1 U
8464 0 0
2
45193.9 0
0
37
1 1 0 0 0 0 0 19 2 0 0 3
347 221
347 425
437 425
2 1 0 0 0 0 0 19 3 0 0 3
365 221
365 383
437 383
3 1 0 0 0 0 0 19 4 0 0 3
401 221
401 340
436 340
4 1 0 0 0 0 0 19 5 0 0 3
419 221
419 298
436 298
5 0 0 0 0 256 0 19 0 0 33 2
374 163
271 163
6 0 0 0 0 256 0 19 0 0 32 3
392 163
392 154
291 154
0 0 1 0 0 4256 0 0 0 0 0 2
712 223
896 223
0 0 1 0 0 32 0 0 0 0 0 2
754 187
754 293
0 0 1 0 0 32 0 0 0 0 0 2
827 187
827 293
0 0 1 0 0 32 0 0 0 0 0 6
717 187
896 187
896 293
712 293
712 187
717 187
0 0 1 0 0 32 0 0 0 0 0 2
732 44
673 44
0 0 1 0 0 32 0 0 0 0 0 2
221 49
300 49
0 0 1 0 0 32 0 0 0 0 0 2
77 49
198 49
0 0 2 0 0 8576 0 0 0 0 0 6
312 132
312 466
693 466
693 106
312 106
312 132
5 0 3 0 0 4096 0 1 0 0 31 2
619 365
682 365
2 0 4 0 0 4096 0 2 0 0 37 2
437 443
130 443
2 0 5 0 0 4096 0 3 0 0 36 2
437 401
150 401
2 0 6 0 0 4096 0 4 0 0 35 2
436 358
170 358
2 0 7 0 0 4096 0 5 0 0 34 2
436 316
190 316
3 3 8 0 0 12416 0 3 1 0 0 4
482 392
524 392
524 370
569 370
3 2 9 0 0 12416 0 4 1 0 0 4
481 349
524 349
524 361
569 361
3 4 10 0 0 8320 0 2 1 0 0 4
482 434
536 434
536 379
569 379
3 1 11 0 0 4224 0 5 1 0 0 4
481 307
536 307
536 352
569 352
2 0 12 0 0 4352 0 9 0 0 33 3
239 113
239 148
271 148
1 0 13 0 0 8448 0 9 0 0 32 3
245 113
245 132
291 132
1 0 4 0 0 0 0 14 0 0 37 3
102 348
102 355
130 355
1 0 5 0 0 0 0 15 0 0 36 3
102 275
102 284
150 284
1 0 6 0 0 0 0 16 0 0 35 3
101 198
101 209
170 209
1 0 7 0 0 0 0 17 0 0 34 3
100 115
100 128
190 128
1 0 3 0 0 0 0 18 0 0 31 3
726 112
726 139
682 139
1 0 3 0 0 4224 0 6 0 0 0 2
682 105
682 613
1 0 13 0 0 4480 0 8 0 0 0 2
291 111
291 612
1 0 12 0 0 4480 0 7 0 0 0 2
271 111
271 612
1 0 7 0 0 4224 0 10 0 0 0 2
190 112
190 612
1 0 6 0 0 4224 0 11 0 0 0 2
170 112
170 612
1 0 5 0 0 4224 0 12 0 0 0 2
150 112
150 613
1 0 4 0 0 4224 0 13 0 0 0 2
130 112
130 614
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
455 81 524 105
461 85 517 101
7 Mux.4x1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
115 27 160 51
121 31 153 47
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
677 21 730 45
683 25 723 41
5 Out's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
240 27 285 51
246 31 278 47
4 Ctrl
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
711 188 756 312
717 192 749 288
22 Dec.

 0
 1
 2
 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 96
758 188 899 312
764 192 892 288
96  Ctrl      Out's
S1  S0       Y
0   0       I0
0   1       I1
1   0       I2
1   1       I3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
