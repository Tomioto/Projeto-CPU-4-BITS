CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
15
12 Hex Display~
7 872 279 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusX
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
9442 0 0
2
45194.8 13
0
14 Logic Display~
6 187 131 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
45194.8 12
0
14 Logic Display~
6 206 131 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
45194.8 11
0
14 Logic Display~
6 226 131 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
45194.8 10
0
14 Logic Display~
6 246 131 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8464 0 0
2
45194.8 9
0
7 Buffer~
58 392 262 0 2 22
0 12 5
0
0 0 96 270
4 4050
-14 -19 14 -11
3 U1D
13 -5 34 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
7168 0 0
2
45194.8 8
0
7 Buffer~
58 445 263 0 2 22
0 11 4
0
0 0 96 270
4 4050
-14 -19 14 -11
3 U1C
13 -5 34 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3171 0 0
2
45194.8 7
0
7 Buffer~
58 496 263 0 2 22
0 10 3
0
0 0 96 270
4 4050
-14 -19 14 -11
3 U1B
13 -5 34 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4139 0 0
2
45194.8 6
0
7 Buffer~
58 549 263 0 2 22
0 9 2
0
0 0 96 270
4 4050
-14 -19 14 -11
3 U1A
13 -5 34 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
6435 0 0
2
45194.8 5
0
14 Logic Display~
6 835 276 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5283 0 0
2
45194.8 4
0
14 Logic Display~
6 815 276 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6874 0 0
2
45194.8 3
0
14 Logic Display~
6 795 276 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5305 0 0
2
45194.8 2
0
14 Logic Display~
6 776 276 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
45194.8 1
0
8 Hex Key~
166 154 124 0 11 12
0 9 10 11 12 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
969 0 0
2
45194.8 0
0
13 MT.Buffer4bit
94 207 267 0 1 17
0 0
13 MT.Buffer4bit
1 0 4736 0
0
2 U2
42 1 56 9
0
0
0
0
0
0
17

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
8402 0 0
2
45193.9 0
0
45
4 0 -1 0 0 16 0 15 0 0 41 2
234 302
234 314
3 0 -1 0 0 16 0 15 0 0 40 2
216 302
216 325
2 0 -1 0 0 16 0 15 0 0 39 2
180 302
180 335
1 0 -1 0 0 16 0 15 0 0 38 2
162 302
162 346
5 0 -1 0 0 16 0 15 0 0 42 2
162 243
162 210
6 0 -1 0 0 16 0 15 0 0 43 2
180 243
180 199
7 0 -1 0 0 16 0 15 0 0 44 2
216 243
216 188
8 0 -1 0 0 16 0 15 0 0 45 2
234 243
234 177
0 0 -1 0 0 48 0 0 0 0 0 2
889 234
767 234
0 0 -1 0 0 48 0 0 0 0 0 2
136 87
254 87
1 0 -1 0 0 16 0 1 0 0 41 2
881 303
881 314
2 0 -1 0 0 16 0 1 0 0 40 2
875 303
875 325
3 0 -1 0 0 16 0 1 0 0 39 2
869 303
869 335
4 0 -1 0 0 16 0 1 0 0 38 2
863 303
863 346
1 0 -1 0 0 16 0 13 0 0 38 2
776 294
776 346
1 0 -1 0 0 16 0 12 0 0 39 2
795 294
795 335
1 0 -1 0 0 16 0 11 0 0 40 2
815 294
815 325
1 0 -1 0 0 16 0 10 0 0 41 2
835 294
835 314
0 0 -1 0 0 272 0 0 0 0 0 5
368 162
368 364
599 364
599 158
368 158
0 0 -1 0 0 272 0 0 0 0 0 5
946 305
980 305
980 359
946 359
946 305
0 0 -1 0 0 272 0 0 0 0 0 5
63 168
97 168
97 222
63 222
63 168
2 0 -1 0 0 16 0 9 0 0 41 2
549 278
549 314
1 0 -1 0 0 16 0 9 0 0 45 2
549 248
549 177
2 0 -1 0 0 16 0 8 0 0 40 2
496 278
496 325
1 0 -1 0 0 16 0 8 0 0 44 2
496 248
496 188
2 0 -1 0 0 16 0 7 0 0 39 2
445 278
445 335
1 0 -1 0 0 16 0 7 0 0 43 2
445 248
445 199
2 0 -1 0 0 16 0 6 0 0 38 2
392 277
392 346
1 0 -1 0 0 16 0 6 0 0 42 2
392 247
392 210
1 0 -1 0 0 16 0 5 0 0 45 2
246 149
246 177
1 0 -1 0 0 16 0 4 0 0 44 2
226 149
226 188
1 0 -1 0 0 16 0 3 0 0 43 2
206 149
206 199
1 0 -1 0 0 16 0 2 0 0 42 2
187 149
187 210
0 0 -1 0 0 16 0 0 0 0 45 2
163 152
163 177
0 0 -1 0 0 16 0 0 0 0 44 2
157 152
157 188
0 0 -1 0 0 16 0 0 0 0 43 2
151 152
151 199
0 0 -1 0 0 16 0 0 0 0 42 2
145 152
145 210
0 0 -1 0 0 16 0 0 0 0 0 2
81 346
967 346
0 0 -1 0 0 16 0 0 0 0 0 2
81 335
967 335
0 0 -1 0 0 16 0 0 0 0 0 2
80 325
966 325
0 0 -1 0 0 16 0 0 0 0 0 2
80 314
966 314
0 0 -1 0 0 16 0 0 0 0 0 2
79 210
614 210
0 0 -1 0 0 16 0 0 0 0 0 2
78 199
614 199
0 0 -1 0 0 16 0 0 0 0 0 2
77 188
614 188
0 0 -1 0 0 16 0 0 0 0 0 2
77 177
614 177
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
442 134 543 158
448 138 536 154
11 Buffer.4bit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
57 147 102 171
63 151 95 167
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
939 284 984 308
945 288 977 304
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
172 62 217 106
178 66 210 98
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
802 210 855 234
808 214 848 230
5 Out's
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
