CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
14
14 Logic Display~
6 120 86 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9265 0 0
2
45194.8 12
0
14 Logic Display~
6 141 86 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9442 0 0
2
45194.8 11
0
14 Logic Display~
6 162 86 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Te
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9424 0 0
2
45194.8 10
0
14 Logic Display~
6 558 86 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 Z
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
45194.8 9
0
14 Logic Display~
6 532 86 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Ts
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9281 0 0
2
45194.8 8
0
9 2-In XOR~
219 317 135 0 3 22
0 5 10 4
0
0 0 96 0
6 74LS86
-21 -24 21 -16
3 U4B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
8464 0 0
2
45194.8 7
0
9 2-In XOR~
219 213 183 0 3 22
0 7 6 10
0
0 0 96 0
6 74LS86
-21 -24 21 -16
3 U4A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
7168 0 0
2
45194.8 6
0
9 2-In AND~
219 326 231 0 3 22
0 10 11 9
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3171 0 0
2
45194.8 5
0
8 2-In OR~
219 429 282 0 3 22
0 9 8 2
0
0 0 96 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
4139 0 0
2
45194.8 4
0
9 Inverter~
13 210 240 0 2 22
0 5 11
0
0 0 96 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
6435 0 0
2
45194.8 3
0
9 2-In AND~
219 219 291 0 3 22
0 6 7 8
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5283 0 0
2
45194.8 2
0
8 Hex Key~
166 68 63 0 11 12
0 7 6 5 14 0 0 0 0 0
4 52
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
6874 0 0
2
45194.8 1
0
12 Hex Display~
7 601 71 0 18 19
10 4 2 12 13 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
5305 0 0
2
45194.8 0
0
10 MT.Sub1bit
94 334 385 0 1 11
0 0
10 MT.Sub1bit
1 0 4736 0
0
2 U5
56 -32 70 -24
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
34 0 0
2
45193.9 0
0
31
2 0 -1 0 0 16 0 14 0 0 28 4
278 386
268 386
268 436
533 436
1 0 -1 0 0 16 0 14 0 0 27 3
334 415
334 422
558 422
3 0 -1 0 0 16 0 14 0 0 29 4
391 385
404 385
404 330
162 330
5 0 -1 0 0 16 0 14 0 0 30 3
357 356
357 346
141 346
4 0 -1 0 0 16 0 14 0 0 31 2
312 357
120 357
3 0 -1 0 0 16 0 9 0 0 28 2
462 282
533 282
0 0 -1 0 0 48 0 0 0 0 0 5
671 311
671 354
917 354
917 311
671 311
0 0 -1 0 0 48 0 0 0 0 0 5
670 138
923 138
923 301
670 301
670 138
0 0 -1 0 0 272 0 0 0 0 0 5
104 104
576 104
576 316
104 316
104 104
0 0 -1 0 0 16 0 0 0 0 28 3
606 107
606 142
533 142
0 0 -1 0 0 16 0 0 0 0 27 3
612 107
612 150
558 150
0 0 -1 0 0 16 0 0 0 0 31 3
66 106
66 159
120 159
0 0 -1 0 0 16 0 0 0 0 30 3
72 106
72 149
141 149
0 0 -1 0 0 16 0 0 0 0 29 3
78 106
78 139
162 139
3 0 -1 0 0 16 0 6 0 0 27 2
350 135
558 135
2 0 -1 0 0 16 0 11 0 0 29 2
195 300
162 300
1 0 -1 0 0 16 0 11 0 0 30 2
195 282
141 282
2 3 -1 0 0 16 0 9 11 0 0 2
416 291
240 291
3 1 -1 0 0 16 0 8 9 0 0 4
347 231
392 231
392 273
416 273
0 1 -1 0 0 272 0 0 8 21 0 3
282 183
282 222
302 222
3 2 -1 0 0 16 0 7 6 0 0 4
246 183
282 183
282 144
301 144
2 2 -1 0 0 16 0 10 8 0 0 2
231 240
302 240
1 0 -1 0 0 16 0 10 0 0 31 2
195 240
120 240
2 0 -1 0 0 16 0 7 0 0 30 2
197 192
141 192
1 0 -1 0 0 16 0 7 0 0 29 2
197 174
162 174
1 0 -1 0 0 16 0 6 0 0 31 2
301 126
120 126
1 0 -1 0 0 16 0 4 0 0 0 2
558 104
558 446
1 0 -1 0 0 16 0 5 0 0 0 4
532 104
532 142
533 142
533 445
1 0 -1 0 0 16 0 3 0 0 0 2
162 104
162 442
1 0 -1 0 0 16 0 2 0 0 0 2
141 104
141 443
1 0 -1 0 0 16 0 1 0 0 0 2
120 104
120 444
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
299 78 368 102
305 82 361 98
7 Sub1bit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 30
882 160 911 324
888 164 904 292
30  0
-1
-1
-2
 1
 0
 0
-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
686 160 707 324
692 164 700 292
22 0
1
2
3
4
5
6
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
673 142 718 166
679 146 711 162
4 Dec.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
878 141 923 165
884 145 916 161
4 Dec.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 49
683 311 912 355
689 315 905 347
49 Z = A (+) (B (+) Te)
Ts = B.Te + ~A . (B (+) Te)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 52
817 143 862 327
823 147 855 291
52 Ts Z
0  0
1  1
1  1
1  0
0  1
0  0
0  0
1  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 63
730 143 791 327
736 147 784 291
63 A B Te
0 0 0 
0 0 1
0 1 0
0 1 1
1 0 0
1 0 1
1 1 0
1 1 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
