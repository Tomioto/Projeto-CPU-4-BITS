CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
22
10 MT.Sub1bit
94 683 414 0 1 11
0 0
10 MT.Sub1bit
9 0 4736 0
0
2 U4
56 -32 70 -24
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
969 0 0
2
45194.8 59
0
10 MT.Sub1bit
94 558 415 0 1 11
0 0
10 MT.Sub1bit
8 0 4736 0
0
2 U3
56 -32 70 -24
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
8402 0 0
2
45194.8 45
0
10 MT.Sub1bit
94 433 416 0 1 11
0 0
10 MT.Sub1bit
7 0 4736 0
0
2 U2
56 -32 70 -24
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
3751 0 0
2
45194.8 31
0
10 MT.Sub1bit
94 307 417 0 1 11
0 0
10 MT.Sub1bit
6 0 4736 0
0
2 U1
56 -32 70 -24
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
4292 0 0
2
45194.8 17
0
12 Hex Display~
7 1016 453 0 16 19
10 2 3 4 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6118 0 0
2
45194.8 16
0
14 Logic Display~
6 173 80 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
34 0 0
2
45194.8 15
0
14 Logic Display~
6 195 80 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6357 0 0
2
45194.8 14
0
14 Logic Display~
6 218 80 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
319 0 0
2
45194.8 13
0
14 Logic Display~
6 239 80 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3976 0 0
2
45194.8 12
0
14 Logic Display~
6 359 78 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7634 0 0
2
45194.8 11
0
14 Logic Display~
6 379 78 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
45194.8 10
0
14 Logic Display~
6 400 78 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6748 0 0
2
45194.8 9
0
14 Logic Display~
6 421 78 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6901 0 0
2
45194.8 8
0
14 Logic Display~
6 958 438 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Z0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
842 0 0
2
45194.8 7
0
14 Logic Display~
6 937 438 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Z1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3277 0 0
2
45194.8 6
0
14 Logic Display~
6 916 438 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Z2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4212 0 0
2
45194.8 5
0
14 Logic Display~
6 896 438 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Z3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4720 0 0
2
45194.8 4
0
7 Ground~
168 763 428 0 1 3
0 0
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5551 0 0
2
45194.8 3
0
14 Logic Display~
6 222 415 0 1 2
10 0
0
0 0 53872 90
6 100MEG
3 -16 45 -8
3 Ts3
-12 -15 9 -7
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6986 0 0
2
45194.8 2
0
8 Hex Key~
166 132 90 0 11 12
0 13 14 15 16 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
8745 0 0
2
45194.8 1
0
8 Hex Key~
166 300 87 0 11 12
0 13 14 15 16 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
9592 0 0
2
45194.8 0
0
10 MT.Sub4bit
94 113 410 0 1 25
0 0
10 MT.Sub4bit
1 0 4736 0
0
2 U5
41 1 55 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
8748 0 0
2
45193.9 0
0
73
4 0 -1 0 0 16 0 22 0 0 47 2
140 445
140 501
3 0 -1 0 0 16 0 22 0 0 45 2
122 445
122 513
2 0 -1 0 0 16 0 22 0 0 46 2
87 445
87 526
1 0 -1 0 0 16 0 22 0 0 44 2
69 445
69 539
9 0 -1 0 0 16 0 22 0 0 70 2
113 386
113 314
10 0 -1 0 0 16 0 22 0 0 71 2
122 386
122 301
11 0 -1 0 0 16 0 22 0 0 72 2
131 386
131 287
12 0 -1 0 0 16 0 22 0 0 73 2
140 386
140 273
5 0 -1 0 0 16 0 22 0 0 66 2
69 386
69 208
6 0 -1 0 0 16 0 22 0 0 67 2
78 386
78 195
7 0 -1 0 0 16 0 22 0 0 68 2
87 386
87 181
8 0 -1 0 0 16 0 22 0 0 69 2
96 386
96 167
1 2 -1 0 0 16 0 19 4 0 0 2
237 418
251 418
1 0 -1 0 0 16 0 1 0 0 47 2
683 444
683 501
1 0 -1 0 0 16 0 2 0 0 45 2
558 445
558 513
1 0 -1 0 0 16 0 3 0 0 46 2
433 446
433 526
1 0 -1 0 0 16 0 4 0 0 44 2
307 447
307 539
5 0 -1 0 0 16 0 1 0 0 73 2
706 385
706 273
4 0 -1 0 0 16 0 1 0 0 69 2
661 386
661 167
5 0 -1 0 0 16 0 2 0 0 72 2
581 386
581 287
4 0 -1 0 0 16 0 2 0 0 68 2
536 387
536 181
5 0 -1 0 0 16 0 3 0 0 71 2
456 387
456 301
4 0 -1 0 0 16 0 3 0 0 67 2
411 388
411 195
5 0 -1 0 0 16 0 4 0 0 70 2
330 388
330 314
4 0 -1 0 0 16 0 4 0 0 66 2
285 389
285 208
3 1 -1 0 0 16 0 1 18 0 0 3
740 414
763 414
763 422
3 2 -1 0 0 16 0 2 1 0 0 2
615 415
627 415
3 2 -1 0 0 16 0 3 2 0 0 2
490 416
502 416
3 2 -1 0 0 16 0 4 3 0 0 2
364 417
377 417
0 0 -1 0 0 48 0 0 0 0 0 2
513 64
770 64
0 0 -1 0 0 48 0 0 0 0 0 2
607 50
607 87
0 0 -1 0 0 48 0 0 0 0 0 5
510 50
770 50
770 87
510 87
510 50
0 0 -1 0 0 48 0 0 0 0 0 2
885 407
1034 407
0 0 -1 0 0 48 0 0 0 0 0 2
115 51
431 51
1 0 -1 0 0 16 0 5 0 0 47 2
1025 477
1025 501
2 0 -1 0 0 16 0 5 0 0 45 2
1019 477
1019 513
3 0 -1 0 0 16 0 5 0 0 46 2
1013 477
1013 526
4 0 -1 0 0 16 0 5 0 0 44 2
1007 477
1007 539
1 0 -1 0 0 16 0 14 0 0 47 2
958 456
958 501
1 0 -1 0 0 16 0 15 0 0 45 2
937 456
937 513
1 0 -1 0 0 16 0 16 0 0 46 2
916 456
916 526
1 0 -1 0 0 16 0 17 0 0 44 2
896 456
896 539
0 0 -1 0 0 272 0 0 0 0 0 6
1053 490
1053 554
1110 554
1110 481
1053 481
1053 490
0 0 -1 0 0 16 0 0 0 0 0 2
28 539
1084 539
0 0 -1 0 0 16 0 0 0 0 0 2
29 513
1085 513
0 0 -1 0 0 16 0 0 0 0 0 2
30 526
1084 526
0 0 -1 0 0 16 0 0 0 0 0 2
29 501
1085 501
0 0 -1 0 0 272 0 0 0 0 0 6
890 264
890 328
947 328
947 255
890 255
890 264
0 0 -1 0 0 272 0 0 0 0 0 6
889 155
889 221
947 221
947 149
889 149
889 155
1 0 -1 0 0 16 0 13 0 0 73 2
421 96
421 273
1 0 -1 0 0 16 0 12 0 0 72 2
400 96
400 287
1 0 -1 0 0 16 0 11 0 0 71 2
379 96
379 301
1 0 -1 0 0 16 0 10 0 0 70 2
359 96
359 314
0 0 -1 0 0 16 0 0 0 0 69 2
309 116
309 167
0 0 -1 0 0 16 0 0 0 0 68 2
303 116
303 181
0 0 -1 0 0 16 0 0 0 0 67 2
297 116
297 195
0 0 -1 0 0 16 0 0 0 0 66 2
291 116
291 208
1 0 -1 0 0 16 0 9 0 0 69 2
239 98
239 167
1 0 -1 0 0 16 0 8 0 0 68 2
218 98
218 181
1 0 -1 0 0 16 0 7 0 0 67 2
195 98
195 195
1 0 -1 0 0 16 0 6 0 0 66 2
173 98
173 208
0 0 -1 0 0 16 0 0 0 0 69 2
141 119
141 167
0 0 -1 0 0 16 0 0 0 0 68 2
135 119
135 181
0 0 -1 0 0 16 0 0 0 0 67 2
129 119
129 195
0 0 -1 0 0 16 0 0 0 0 66 2
123 119
123 208
0 0 -1 0 0 16 0 0 0 0 0 2
26 208
909 208
0 0 -1 0 0 16 0 0 0 0 0 2
27 195
909 195
0 0 -1 0 0 16 0 0 0 0 0 2
27 181
910 181
0 0 -1 0 0 16 0 0 0 0 0 2
25 167
911 167
0 0 -1 0 0 16 0 0 0 0 0 2
27 314
910 314
0 0 -1 0 0 16 0 0 0 0 0 2
28 301
910 301
0 0 -1 0 0 16 0 0 0 0 0 2
28 287
911 287
0 0 -1 0 0 16 0 0 0 0 0 2
26 273
912 273
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
888 126 933 150
894 130 926 146
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
238 27 283 51
244 31 276 47
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
932 383 985 407
938 387 978 403
5 Out's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1052 458 1097 482
1058 462 1090 478
4 BusZ
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
889 233 934 257
895 237 927 253
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 58
503 46 772 90
509 50 765 82
58    In's            Out's
 BusA, BusB   Busz = BusA + BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
511 113 700 137
517 117 693 133
22 * Subtrator Aritm�tico
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
578 25 663 49
584 29 656 45
9 Sub.4bits
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
