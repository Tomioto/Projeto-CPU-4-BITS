CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
8388626 0
0
6 Title:
5 Name:
0
0
0
13
9 2-In AND~
219 257 314 0 3 22
0 6 7 8
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
3284 0 0
2
45189.9 0
0
9 Inverter~
13 248 263 0 2 22
0 5 11
0
0 0 112 0
6 74LS04
-21 -19 21 -11
3 U4A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 4 0
1 U
659 0 0
2
45189.9 0
0
8 2-In OR~
219 467 305 0 3 22
0 9 8 2
0
0 0 112 0
6 74LS32
-21 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3800 0 0
2
45189.9 0
0
9 2-In AND~
219 364 254 0 3 22
0 10 11 9
0
0 0 112 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6792 0 0
2
45189.9 0
0
9 2-In XOR~
219 251 206 0 3 22
0 7 6 10
0
0 0 112 0
6 74LS86
-21 -24 21 -16
3 U1B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3701 0 0
2
45189.9 0
0
9 2-In XOR~
219 355 158 0 3 22
0 5 10 4
0
0 0 112 0
6 74LS86
-21 -24 21 -16
3 U1A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6316 0 0
2
45189.9 0
0
14 Logic Display~
6 570 109 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Ts
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8734 0 0
2
45189.9 0
0
14 Logic Display~
6 596 109 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 Z
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7988 0 0
2
45189.9 0
0
14 Logic Display~
6 200 109 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Te
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3217 0 0
2
45189.9 0
0
14 Logic Display~
6 179 109 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3965 0 0
2
45189.9 0
0
14 Logic Display~
6 158 109 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8239 0 0
2
45189.9 0
0
12 Hex Display~
7 641 106 0 18 19
10 4 2 12 13 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
828 0 0
2
45189.9 0
0
8 Hex Key~
166 107 105 0 11 12
0 7 6 5 14 0 0 0 0 0
4 52
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
3 KPD
6187 0 0
2
45189.9 0
0
26
3 0 2 0 0 4096 0 3 0 0 23 2
500 305
571 305
0 0 1 0 0 8224 0 0 0 0 0 5
709 334
709 377
955 377
955 334
709 334
0 0 1 0 0 4256 0 0 0 0 0 5
708 161
961 161
961 324
708 324
708 161
0 0 3 0 0 4480 0 0 0 0 0 5
142 127
614 127
614 339
142 339
142 127
2 0 2 0 0 8192 0 12 0 0 23 3
644 130
644 165
571 165
1 0 4 0 0 8192 0 12 0 0 22 3
650 130
650 173
596 173
3 0 5 0 0 8192 0 13 0 0 26 3
104 129
104 182
158 182
2 0 6 0 0 8192 0 13 0 0 25 3
110 129
110 172
179 172
1 0 7 0 0 8192 0 13 0 0 24 3
116 129
116 162
200 162
3 0 4 0 0 4096 0 6 0 0 22 2
388 158
596 158
2 0 7 0 0 0 0 1 0 0 24 2
233 323
200 323
1 0 6 0 0 0 0 1 0 0 25 2
233 305
179 305
2 3 8 0 0 4224 0 3 1 0 0 2
454 314
278 314
3 1 9 0 0 4224 0 4 3 0 0 4
385 254
430 254
430 296
454 296
0 1 10 0 0 4480 0 0 4 16 0 3
320 206
320 245
340 245
3 2 10 0 0 0 0 5 6 0 0 4
284 206
320 206
320 167
339 167
2 2 11 0 0 4224 0 2 4 0 0 2
269 263
340 263
1 0 5 0 0 4096 0 2 0 0 26 2
233 263
158 263
2 0 6 0 0 0 0 5 0 0 25 2
235 215
179 215
1 0 7 0 0 0 0 5 0 0 24 2
235 197
200 197
1 0 5 0 0 4096 0 6 0 0 26 2
339 149
158 149
1 0 4 0 0 4224 0 8 0 0 0 2
596 127
596 469
1 0 2 0 0 12416 0 7 0 0 0 4
570 127
570 165
571 165
571 468
1 0 7 0 0 4224 0 9 0 0 0 2
200 127
200 465
1 0 6 0 0 4224 0 10 0 0 0 2
179 127
179 466
1 0 5 0 0 4224 0 11 0 0 0 2
158 127
158 467
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 30
920 183 949 347
926 187 942 315
30  0
-1
-1
-2
 1
 0
 0
-1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
724 183 745 347
730 187 738 315
22 0
1
2
3
4
5
6
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
711 165 756 189
717 169 749 185
4 Dec.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
916 164 961 188
922 168 954 184
4 Dec.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 49
721 334 950 378
727 338 943 370
49 Z = A (+) (B (+) Te)
Ts = B.Te + ~A . (B (+) Te)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 52
855 166 900 350
861 170 893 314
52 Ts Z
0  0
1  1
1  1
1  0
0  1
0  0
0  0
1  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 63
768 166 829 350
774 170 822 314
63 A B Te
0 0 0 
0 0 1
0 1 0
0 1 1
1 0 0
1 0 1
1 1 0
1 1 1
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
