CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
27
9 MT.Mux4x1
94 573 562 0 7 15
0 15 18 21 26 5 10 9
9 MT.Mux4x1
17 0 4224 0
0
2 U8
50 0 64 8
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
7168 0 0
2
45194.8 299
0
9 MT.Mux4x1
94 430 565 0 7 15
0 16 19 22 25 6 10 9
9 MT.Mux4x1
16 0 4224 0
0
2 U7
50 0 64 8
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
631 0 0
2
45194.8 265
0
9 MT.Mux4x1
94 295 565 0 7 15
0 17 20 23 24 7 10 9
9 MT.Mux4x1
15 0 4224 0
0
2 U6
50 0 64 8
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
9466 0 0
2
45194.8 231
0
9 MT.Mux4x1
94 152 567 0 7 15
0 12 11 13 14 8 10 9
9 MT.Mux4x1
14 0 4224 0
0
2 U5
50 0 64 8
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3266 0 0
2
45194.8 197
0
10 MT.Add4bit
94 529 257 0 12 25
0 14 24 25 26 31 32 33 34 27
28 29 30
10 MT.Add4bit
13 0 4224 0
0
2 U4
42 0 56 8
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
7693 0 0
2
45194.8 127
0
13 MT.Buffer4bit
94 407 256 0 8 17
0 13 23 22 21 31 32 33 34
13 MT.Buffer4bit
12 0 4224 0
0
2 U3
42 1 56 9
0
0
0
0
0
0
17

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3723 0 0
2
45194.8 112
0
12 MT.Nand4bits
94 286 256 0 12 25
0 11 20 19 18 31 32 33 34 27
28 29 30
12 MT.Nand4bits
11 0 4224 0
0
2 U2
42 1 56 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3440 0 0
2
45194.8 92
0
10 MT.Sub4bit
94 165 254 0 12 25
0 12 17 16 15 31 32 33 34 27
28 29 30
10 MT.Sub4bit
10 0 4224 0
0
2 U1
41 1 55 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
6263 0 0
2
45194.8 18
0
8 Hex Key~
166 564 80 0 11 12
0 34 33 32 31 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
4900 0 0
2
45194.8 17
0
8 Hex Key~
166 718 81 0 11 12
0 172 29 28 27 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
8783 0 0
2
45194.8 16
0
14 Logic Display~
6 599 82 0 1 2
10 31
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3221 0 0
2
45194.8 15
0
14 Logic Display~
6 619 82 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3215 0 0
2
45194.8 14
0
14 Logic Display~
6 639 82 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7903 0 0
2
45194.8 13
0
14 Logic Display~
6 659 82 0 1 2
10 34
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7121 0 0
2
45194.8 12
0
14 Logic Display~
6 815 81 0 1 2
10 30
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4484 0 0
2
45194.8 11
0
14 Logic Display~
6 755 81 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5996 0 0
2
45194.8 10
0
14 Logic Display~
6 775 81 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7804 0 0
2
45194.8 9
0
14 Logic Display~
6 795 81 0 1 2
10 29
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5523 0 0
2
45194.8 8
0
12 Hex Display~
7 873 619 0 16 19
10 5 6 7 8 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3330 0 0
2
45194.8 7
0
14 Logic Display~
6 948 623 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3465 0 0
2
45194.8 6
0
14 Logic Display~
6 928 623 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8396 0 0
2
45194.8 5
0
14 Logic Display~
6 908 623 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3685 0 0
2
45194.8 4
0
14 Logic Display~
6 968 623 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7849 0 0
2
45194.8 3
0
8 Hex Key~
166 720 587 0 11 12
0 10 9 170 171 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
6343 0 0
2
45194.8 2
0
14 Logic Display~
6 771 593 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7376 0 0
2
45194.8 1
0
14 Logic Display~
6 751 593 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9156 0 0
2
45194.8 0
0
10 MT.ULA4bit
94 644 254 0 1 29
0 0
10 MT.ULA4bit
1 0 4736 0
0
2 U9
-89 3 -75 11
0
0
0
0
0
0
29

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
5776 0 0
2
45194.1 0
0
157
5 0 -1 0 0 272 0 27 0 0 125 6
695 271
695 270
789 270
789 659
677 659
677 638
6 0 -1 0 0 272 0 27 0 0 124 6
704 254
704 253
802 253
802 650
694 650
694 622
0 0 -1 0 0 48 0 0 0 0 0 2
837 318
1080 318
0 0 -1 0 0 48 0 0 0 0 0 2
950 298
950 389
0 0 -1 0 0 48 0 0 0 0 0 2
879 298
879 389
0 0 -1 0 0 48 0 0 0 0 0 5
837 298
1080 298
1080 389
837 389
837 298
4 0 -1 0 0 16 0 27 0 0 149 2
653 295
653 666
3 0 -1 0 0 16 0 27 0 0 148 2
644 295
644 676
2 0 -1 0 0 16 0 27 0 0 147 2
635 295
635 687
1 0 -1 0 0 16 0 27 0 0 146 2
626 295
626 698
11 0 -1 0 0 16 0 27 0 0 150 2
671 228
671 192
12 0 -1 0 0 16 0 27 0 0 151 2
680 228
680 183
13 0 -1 0 0 16 0 27 0 0 152 2
689 228
689 174
14 0 -1 0 0 16 0 27 0 0 153 2
698 228
698 165
7 0 -1 0 0 16 0 27 0 0 154 4
583 228
583 221
577 221
577 145
8 0 -1 0 0 16 0 27 0 0 155 4
593 228
593 216
586 216
586 136
9 0 -1 0 0 16 0 27 0 0 156 4
601 228
601 205
593 205
593 127
10 0 -1 0 0 16 0 27 0 0 157 2
610 228
610 118
0 0 -1 0 0 48 0 0 0 0 0 2
549 36
825 36
0 0 -1 0 0 48 0 0 0 0 0 2
850 573
985 573
0 0 -1 0 0 48 0 0 0 0 0 2
705 545
783 545
0 0 -1 0 0 272 0 0 0 0 0 5
823 159
823 204
862 204
862 159
823 159
0 0 -1 0 0 272 0 0 0 0 0 5
981 657
981 710
1018 710
1018 657
981 657
1 0 -1 0 0 16 0 23 0 0 149 2
968 641
968 666
1 0 -1 0 0 16 0 20 0 0 148 2
948 641
948 676
1 0 -1 0 0 16 0 21 0 0 147 2
928 641
928 687
1 0 -1 0 0 16 0 22 0 0 146 2
908 641
908 698
1 0 -1 0 0 16 0 19 0 0 149 2
882 643
882 666
2 0 -1 0 0 16 0 19 0 0 148 2
876 643
876 676
3 0 -1 0 0 16 0 19 0 0 147 2
870 643
870 687
4 0 -1 0 0 16 0 19 0 0 146 2
864 643
864 698
1 0 -1 0 0 272 0 26 0 0 125 2
751 611
751 638
1 0 -1 0 0 272 0 25 0 0 124 2
771 611
771 622
2 0 -1 0 0 272 0 24 0 0 125 2
723 611
723 638
1 0 -1 0 0 272 0 24 0 0 124 2
729 611
729 622
5 0 -1 0 0 16 0 1 0 0 149 2
573 596
573 666
5 0 -1 0 0 16 0 2 0 0 148 2
430 599
430 676
5 0 -1 0 0 16 0 3 0 0 147 2
295 599
295 687
5 0 -1 0 0 16 0 4 0 0 146 2
152 601
152 698
7 0 -1 0 0 272 0 1 0 0 125 2
521 571
521 638
6 0 -1 0 0 272 0 1 0 0 124 3
521 562
501 562
501 622
7 0 -1 0 0 272 0 2 0 0 125 2
378 574
378 638
6 0 -1 0 0 272 0 2 0 0 124 3
378 565
356 565
356 622
7 0 -1 0 0 272 0 3 0 0 125 3
243 574
230 574
230 638
6 0 -1 0 0 272 0 3 0 0 124 3
243 565
216 565
216 622
7 0 -1 0 0 272 0 4 0 0 125 2
100 576
100 638
6 0 -1 0 0 272 0 4 0 0 124 3
100 567
86 567
86 622
2 0 -1 0 0 16 0 4 0 0 134 4
134 542
134 529
129 529
129 455
1 0 -1 0 0 16 0 4 0 0 138 4
116 542
116 530
109 530
109 506
3 0 -1 0 0 16 0 4 0 0 142 4
170 542
170 529
162 529
162 401
4 0 -1 0 0 16 0 4 0 0 130 4
188 542
188 522
182 522
182 347
4 0 -1 0 0 16 0 8 0 0 141 2
192 289
192 476
3 0 -1 0 0 16 0 8 0 0 140 2
174 289
174 486
2 0 -1 0 0 16 0 8 0 0 139 2
139 289
139 496
1 0 -1 0 0 16 0 8 0 0 138 2
121 289
121 506
4 0 -1 0 0 16 0 7 0 0 137 4
313 291
313 305
306 305
306 425
3 0 -1 0 0 16 0 7 0 0 136 2
295 291
295 435
2 0 -1 0 0 16 0 7 0 0 135 2
259 291
259 445
1 0 -1 0 0 16 0 7 0 0 134 2
242 291
242 455
4 0 -1 0 0 16 0 6 0 0 145 2
434 291
434 371
3 0 -1 0 0 16 0 6 0 0 144 2
416 291
416 381
2 0 -1 0 0 16 0 6 0 0 143 2
380 291
380 391
1 0 -1 0 0 16 0 6 0 0 142 2
362 291
362 401
1 0 -1 0 0 16 0 3 0 0 139 2
259 540
259 496
2 0 -1 0 0 16 0 3 0 0 135 2
277 540
277 445
3 0 -1 0 0 16 0 3 0 0 143 2
313 540
313 391
4 0 -1 0 0 16 0 3 0 0 131 2
331 540
331 337
1 0 -1 0 0 16 0 2 0 0 140 2
394 540
394 486
2 0 -1 0 0 16 0 2 0 0 136 2
412 540
412 435
3 0 -1 0 0 16 0 2 0 0 144 2
448 540
448 381
4 0 -1 0 0 16 0 2 0 0 132 2
466 540
466 327
1 0 -1 0 0 16 0 1 0 0 141 2
537 537
537 476
2 0 -1 0 0 16 0 1 0 0 137 2
555 537
555 425
3 0 -1 0 0 16 0 1 0 0 145 2
591 537
591 371
4 0 -1 0 0 16 0 1 0 0 133 2
609 537
609 317
4 0 -1 0 0 16 0 5 0 0 133 2
556 290
556 317
3 0 -1 0 0 16 0 5 0 0 132 2
538 290
538 327
2 0 -1 0 0 16 0 5 0 0 131 2
502 290
502 337
1 0 -1 0 0 16 0 5 0 0 130 2
484 290
484 347
9 0 -1 0 0 16 0 5 0 0 150 2
529 233
529 192
10 0 -1 0 0 16 0 5 0 0 151 2
538 233
538 183
11 0 -1 0 0 16 0 5 0 0 152 2
547 233
547 174
12 0 -1 0 0 16 0 5 0 0 153 2
557 233
557 165
5 0 -1 0 0 16 0 5 0 0 154 2
484 233
484 145
6 0 -1 0 0 16 0 5 0 0 155 2
493 233
493 136
7 0 -1 0 0 16 0 5 0 0 156 2
503 233
503 127
8 0 -1 0 0 16 0 5 0 0 157 2
512 233
512 118
5 0 -1 0 0 16 0 6 0 0 154 2
362 232
362 145
6 0 -1 0 0 16 0 6 0 0 155 2
380 232
380 136
7 0 -1 0 0 16 0 6 0 0 156 2
416 232
416 127
8 0 -1 0 0 16 0 6 0 0 157 2
434 232
434 118
9 0 -1 0 0 16 0 7 0 0 150 2
286 232
286 192
10 0 -1 0 0 16 0 7 0 0 151 2
295 232
295 183
11 0 -1 0 0 16 0 7 0 0 152 2
304 232
304 174
12 0 -1 0 0 16 0 7 0 0 153 2
313 232
313 165
5 0 -1 0 0 16 0 7 0 0 154 2
241 232
241 145
6 0 -1 0 0 16 0 7 0 0 155 2
251 232
251 136
7 0 -1 0 0 16 0 7 0 0 156 2
260 232
260 127
8 0 -1 0 0 16 0 7 0 0 157 2
269 232
269 118
9 0 -1 0 0 16 0 8 0 0 150 2
165 230
165 192
10 0 -1 0 0 16 0 8 0 0 151 2
174 230
174 183
11 0 -1 0 0 16 0 8 0 0 152 2
183 230
183 174
12 0 -1 0 0 16 0 8 0 0 153 2
192 230
192 165
5 0 -1 0 0 16 0 8 0 0 154 2
121 230
121 145
6 0 -1 0 0 16 0 8 0 0 155 2
130 230
130 136
7 0 -1 0 0 16 0 8 0 0 156 2
139 230
139 127
8 0 -1 0 0 16 0 8 0 0 157 2
148 230
148 118
1 0 -1 0 0 16 0 15 0 0 153 2
815 99
815 165
1 0 -1 0 0 16 0 18 0 0 152 2
795 99
795 174
1 0 -1 0 0 16 0 17 0 0 151 2
775 99
775 183
1 0 -1 0 0 16 0 16 0 0 150 2
755 99
755 192
2 0 -1 0 0 16 0 10 0 0 152 2
721 105
721 174
3 0 -1 0 0 16 0 10 0 0 151 2
715 105
715 183
4 0 -1 0 0 16 0 10 0 0 150 4
709 105
709 187
710 187
710 192
1 0 -1 0 0 16 0 14 0 0 157 2
659 100
659 118
1 0 -1 0 0 16 0 13 0 0 156 2
639 100
639 127
1 0 -1 0 0 16 0 12 0 0 155 2
619 100
619 136
1 0 -1 0 0 16 0 11 0 0 154 2
599 100
599 145
1 0 -1 0 0 16 0 9 0 0 157 2
573 104
573 118
2 0 -1 0 0 16 0 9 0 0 156 2
567 104
567 127
3 0 -1 0 0 16 0 9 0 0 155 2
561 104
561 136
4 0 -1 0 0 16 0 9 0 0 154 2
555 104
555 145
0 0 -1 0 0 272 0 0 0 0 0 5
824 112
824 152
861 152
861 108
823 108
0 0 -1 0 0 272 0 0 0 0 0 2
62 622
776 622
0 0 -1 0 0 272 0 0 0 0 0 2
62 638
775 638
0 0 -1 0 0 272 0 0 0 0 0 5
661 470
699 470
699 514
661 514
661 470
0 0 -1 0 0 272 0 0 0 0 0 5
662 420
662 463
699 463
699 416
661 416
0 0 -1 0 0 272 0 0 0 0 0 5
662 364
699 364
699 408
662 408
662 364
0 0 -1 0 0 272 0 0 0 0 0 5
662 304
662 355
698 355
698 304
662 304
0 0 -1 0 0 16 0 0 0 0 0 2
87 347
672 347
0 0 -1 0 0 16 0 0 0 0 0 2
88 337
673 337
0 0 -1 0 0 16 0 0 0 0 0 2
87 327
672 327
0 0 -1 0 0 16 0 0 0 0 0 2
86 317
671 317
0 0 -1 0 0 16 0 0 0 0 0 2
88 455
673 455
0 0 -1 0 0 16 0 0 0 0 0 2
89 445
674 445
0 0 -1 0 0 16 0 0 0 0 0 2
88 435
673 435
0 0 -1 0 0 16 0 0 0 0 0 2
87 425
672 425
0 0 -1 0 0 16 0 0 0 0 0 2
90 506
675 506
0 0 -1 0 0 16 0 0 0 0 0 2
91 496
676 496
0 0 -1 0 0 16 0 0 0 0 0 2
90 486
675 486
0 0 -1 0 0 16 0 0 0 0 0 2
89 476
674 476
0 0 -1 0 0 16 0 0 0 0 0 2
90 401
675 401
0 0 -1 0 0 16 0 0 0 0 0 2
91 391
676 391
0 0 -1 0 0 16 0 0 0 0 0 2
90 381
675 381
0 0 -1 0 0 16 0 0 0 0 0 2
89 371
674 371
0 0 -1 0 0 16 0 0 0 0 0 2
17 698
990 698
0 0 -1 0 0 16 0 0 0 0 0 2
17 687
991 687
0 0 -1 0 0 16 0 0 0 0 0 2
17 676
990 676
0 0 -1 0 0 16 0 0 0 0 0 2
17 666
991 666
0 0 -1 0 0 16 0 0 0 0 0 2
18 192
839 192
0 0 -1 0 0 16 0 0 0 0 0 2
17 183
839 183
0 0 -1 0 0 16 0 0 0 0 0 2
18 174
839 174
0 0 -1 0 0 16 0 0 0 0 0 2
18 165
840 165
0 0 -1 0 0 16 0 0 0 0 0 2
16 145
837 145
0 0 -1 0 0 16 0 0 0 0 0 2
15 136
837 136
0 0 -1 0 0 16 0 0 0 0 0 2
16 127
837 127
0 0 -1 0 0 16 0 0 0 0 0 2
16 118
838 118
18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
982 255 1047 299
986 259 1042 291
14 Funcoes
Out`s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
893 256 934 300
897 260 929 292
10 Ctrl
In`s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 98
881 299 1082 403
885 303 1077 383
98 S1  S0    BusU
 0   0    BusA+BusB
 0   1    BusA
 1   0    BusA.BusB(neg)
 1   1    BusA-BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
838 298 879 402
842 302 874 382
20 Dec.
 0
 1
 2
 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
699 302 740 326
703 306 735 322
4 BusW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
701 362 742 386
705 366 737 382
4 BusX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
701 413 742 437
705 417 737 433
4 BusY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
701 466 742 490
705 470 737 486
4 BusZ
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
701 322 734 346
705 326 729 342
3 Add
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
698 382 755 406
702 386 750 402
6 Buffer
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
701 433 742 457
705 437 737 453
4 Nand
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
701 483 734 507
705 487 729 503
3 Sub
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1020 676 1061 700
1024 680 1056 696
4 BusU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
861 122 902 146
865 126 897 142
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
862 172 903 196
866 176 898 192
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
666 13 707 37
670 17 702 33
4 In`s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
710 525 775 549
714 529 770 545
7 Funcoes
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
893 551 942 575
897 555 937 571
5 Out`s
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
