CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
8388626 0
0
6 Title:
5 Name:
0
0
0
26
14 Logic Display~
6 748 611 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.90094e-315 5.26354e-315
0
14 Logic Display~
6 768 611 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.90094e-315 0
0
8 Hex Key~
166 717 605 0 11 12
0 10 9 170 171 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD3
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
7361 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 965 641 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.90094e-315 5.32571e-315
0
14 Logic Display~
6 905 641 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90094e-315 5.30499e-315
0
14 Logic Display~
6 925 641 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.90094e-315 5.26354e-315
0
14 Logic Display~
6 945 641 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.90094e-315 0
0
12 Hex Display~
7 870 637 0 16 19
10 5 6 7 8 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3536 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 792 99 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.90094e-315 5.32571e-315
0
14 Logic Display~
6 772 99 0 1 2
10 28
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.90094e-315 5.30499e-315
0
14 Logic Display~
6 752 99 0 1 2
10 27
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90094e-315 5.26354e-315
0
14 Logic Display~
6 812 99 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 656 100 0 1 2
10 34
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 636 100 0 1 2
10 33
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 616 100 0 1 2
10 32
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3108 0 0
2
5.90094e-315 0
0
14 Logic Display~
6 596 100 0 1 2
10 31
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4299 0 0
2
5.90094e-315 0
0
8 Hex Key~
166 715 99 0 11 12
0 172 29 28 27 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD2
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9672 0 0
2
5.90094e-315 0
0
8 Hex Key~
166 561 98 0 11 12
0 34 33 32 31 0 0 0 0 0
0 48
0
0 0 4656 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 1 0 0 0
3 KPD
7876 0 0
2
5.90094e-315 0
0
10 MT.Sub4bit
94 162 272 0 12 25
0 12 17 16 15 31 32 33 34 27
28 29 30
10 MT.Sub4bit
1 0 4240 0
0
2 U1
41 1 55 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
6369 0 0
2
5.90094e-315 0
0
12 MT.Nand4bits
94 283 274 0 12 25
0 11 20 19 18 31 32 33 34 27
28 29 30
12 MT.Nand4bits
2 0 4240 0
0
2 U2
42 1 56 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
9172 0 0
2
5.90094e-315 0
0
13 MT.Buffer4bit
94 404 274 0 8 17
0 13 23 22 21 31 32 33 34
13 MT.Buffer4bit
3 0 4240 0
0
2 U3
42 1 56 9
0
0
0
0
0
0
17

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
7100 0 0
2
5.90094e-315 0
0
10 MT.Add4bit
94 526 275 0 12 25
0 14 24 25 26 31 32 33 34 27
28 29 30
10 MT.Add4bit
4 0 4240 0
0
2 U4
42 0 56 8
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3820 0 0
2
5.90094e-315 0
0
9 MT.Mux4x1
94 149 585 0 7 15
0 12 11 13 14 8 10 9
9 MT.Mux4x1
5 0 4240 0
0
2 U5
50 0 64 8
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
7678 0 0
2
5.90094e-315 0
0
9 MT.Mux4x1
94 292 583 0 7 15
0 17 20 23 24 7 10 9
9 MT.Mux4x1
6 0 4240 0
0
2 U6
50 0 64 8
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
961 0 0
2
5.90094e-315 0
0
9 MT.Mux4x1
94 427 583 0 7 15
0 16 19 22 25 6 10 9
9 MT.Mux4x1
7 0 4240 0
0
2 U7
50 0 64 8
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3178 0 0
2
5.90094e-315 0
0
9 MT.Mux4x1
94 570 580 0 7 15
0 15 18 21 26 5 10 9
9 MT.Mux4x1
8 0 4240 0
0
2 U8
50 0 64 8
0
0
0
0
0
0
15

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 1 0 0 0
1 U
3409 0 0
2
5.90094e-315 0
0
144
1 0 0 0 0 0 0 17 0 0 140 2
724 123
724 183
0 0 1 0 0 4128 0 0 0 0 0 2
755 346
998 346
0 0 1 0 0 32 0 0 0 0 0 2
868 326
868 417
0 0 1 0 0 32 0 0 0 0 0 2
797 326
797 417
0 0 1 0 0 32 0 0 0 0 0 5
755 326
998 326
998 417
755 417
755 326
0 0 1 0 0 4256 0 0 0 0 0 2
546 54
822 54
0 0 1 0 0 32 0 0 0 0 0 2
847 591
982 591
0 0 1 0 0 32 0 0 0 0 0 2
702 563
780 563
0 0 3 0 0 4480 0 0 0 0 0 5
820 177
820 222
859 222
859 177
820 177
0 0 4 0 0 4480 0 0 0 0 0 5
978 675
978 728
1015 728
1015 675
978 675
1 0 5 0 0 4096 0 4 0 0 136 2
965 659
965 684
1 0 6 0 0 4096 0 7 0 0 135 2
945 659
945 694
1 0 7 0 0 4096 0 6 0 0 134 2
925 659
925 705
1 0 8 0 0 4096 0 5 0 0 133 2
905 659
905 716
1 0 5 0 0 0 0 8 0 0 136 2
879 661
879 684
2 0 6 0 0 0 0 8 0 0 135 2
873 661
873 694
3 0 7 0 0 0 0 8 0 0 134 2
867 661
867 705
4 0 8 0 0 0 0 8 0 0 133 2
861 661
861 716
1 0 9 0 0 4352 0 1 0 0 112 2
748 629
748 656
1 0 10 0 0 4352 0 2 0 0 111 2
768 629
768 640
2 0 9 0 0 256 0 3 0 0 112 2
720 629
720 656
1 0 10 0 0 256 0 3 0 0 111 2
726 629
726 640
5 0 5 0 0 4096 0 26 0 0 136 2
570 614
570 684
5 0 6 0 0 4096 0 25 0 0 135 2
427 617
427 694
5 0 7 0 0 4096 0 24 0 0 134 2
292 617
292 705
5 0 8 0 0 4096 0 23 0 0 133 2
149 619
149 716
7 0 9 0 0 4352 0 26 0 0 112 2
518 589
518 656
6 0 10 0 0 8448 0 26 0 0 111 3
518 580
498 580
498 640
7 0 9 0 0 256 0 25 0 0 112 2
375 592
375 656
6 0 10 0 0 256 0 25 0 0 111 3
375 583
353 583
353 640
7 0 9 0 0 256 0 24 0 0 112 3
240 592
227 592
227 656
6 0 10 0 0 256 0 24 0 0 111 3
240 583
213 583
213 640
7 0 9 0 0 256 0 23 0 0 112 2
97 594
97 656
6 0 10 0 0 256 0 23 0 0 111 3
97 585
83 585
83 640
2 0 11 0 0 12288 0 23 0 0 121 4
131 560
131 547
126 547
126 473
1 0 12 0 0 12288 0 23 0 0 125 4
113 560
113 548
106 548
106 524
3 0 13 0 0 12288 0 23 0 0 129 4
167 560
167 547
159 547
159 419
4 0 14 0 0 12288 0 23 0 0 117 4
185 560
185 540
179 540
179 365
4 0 15 0 0 4096 0 19 0 0 128 2
189 307
189 494
3 0 16 0 0 4096 0 19 0 0 127 2
171 307
171 504
2 0 17 0 0 4096 0 19 0 0 126 2
136 307
136 514
1 0 12 0 0 4096 0 19 0 0 125 2
118 307
118 524
4 0 18 0 0 12288 0 20 0 0 124 4
310 309
310 323
303 323
303 443
3 0 19 0 0 4096 0 20 0 0 123 2
292 309
292 453
2 0 20 0 0 4096 0 20 0 0 122 2
256 309
256 463
1 0 11 0 0 4096 0 20 0 0 121 2
239 309
239 473
4 0 21 0 0 4096 0 21 0 0 132 2
431 309
431 389
3 0 22 0 0 4096 0 21 0 0 131 2
413 309
413 399
2 0 23 0 0 4096 0 21 0 0 130 2
377 309
377 409
1 0 13 0 0 0 0 21 0 0 129 2
359 309
359 419
1 0 17 0 0 0 0 24 0 0 126 2
256 558
256 514
2 0 20 0 0 0 0 24 0 0 122 2
274 558
274 463
3 0 23 0 0 4096 0 24 0 0 130 2
310 558
310 409
4 0 24 0 0 4096 0 24 0 0 118 2
328 558
328 355
1 0 16 0 0 0 0 25 0 0 127 2
391 558
391 504
2 0 19 0 0 0 0 25 0 0 123 2
409 558
409 453
3 0 22 0 0 4096 0 25 0 0 131 2
445 558
445 399
4 0 25 0 0 4096 0 25 0 0 119 2
463 558
463 345
1 0 15 0 0 0 0 26 0 0 128 2
534 555
534 494
2 0 18 0 0 0 0 26 0 0 124 2
552 555
552 443
3 0 21 0 0 4096 0 26 0 0 132 2
588 555
588 389
4 0 26 0 0 4096 0 26 0 0 120 2
606 555
606 335
4 0 26 0 0 0 0 22 0 0 120 2
553 308
553 335
3 0 25 0 0 0 0 22 0 0 119 2
535 308
535 345
2 0 24 0 0 0 0 22 0 0 118 2
499 308
499 355
1 0 14 0 0 0 0 22 0 0 117 2
481 308
481 365
9 0 27 0 0 4096 0 22 0 0 137 2
526 251
526 210
10 0 28 0 0 4096 0 22 0 0 138 2
535 251
535 201
11 0 29 0 0 4096 0 22 0 0 139 2
544 251
544 192
12 0 30 0 0 4096 0 22 0 0 140 2
554 251
554 183
5 0 31 0 0 4096 0 22 0 0 141 2
481 251
481 163
6 0 32 0 0 4096 0 22 0 0 142 2
490 251
490 154
7 0 33 0 0 4096 0 22 0 0 143 2
500 251
500 145
8 0 34 0 0 4096 0 22 0 0 144 2
509 251
509 136
5 0 31 0 0 0 0 21 0 0 141 2
359 250
359 163
6 0 32 0 0 0 0 21 0 0 142 2
377 250
377 154
7 0 33 0 0 0 0 21 0 0 143 2
413 250
413 145
8 0 34 0 0 0 0 21 0 0 144 2
431 250
431 136
9 0 27 0 0 0 0 20 0 0 137 2
283 250
283 210
10 0 28 0 0 0 0 20 0 0 138 2
292 250
292 201
11 0 29 0 0 0 0 20 0 0 139 2
301 250
301 192
12 0 30 0 0 0 0 20 0 0 140 2
310 250
310 183
5 0 31 0 0 0 0 20 0 0 141 2
238 250
238 163
6 0 32 0 0 0 0 20 0 0 142 2
248 250
248 154
7 0 33 0 0 0 0 20 0 0 143 2
257 250
257 145
8 0 34 0 0 0 0 20 0 0 144 2
266 250
266 136
9 0 27 0 0 0 0 19 0 0 137 2
162 248
162 210
10 0 28 0 0 0 0 19 0 0 138 2
171 248
171 201
11 0 29 0 0 0 0 19 0 0 139 2
180 248
180 192
12 0 30 0 0 0 0 19 0 0 140 2
189 248
189 183
5 0 31 0 0 0 0 19 0 0 141 2
118 248
118 163
6 0 32 0 0 0 0 19 0 0 142 2
127 248
127 154
7 0 33 0 0 0 0 19 0 0 143 2
136 248
136 145
8 0 34 0 0 0 0 19 0 0 144 2
145 248
145 136
1 0 30 0 0 0 0 12 0 0 140 2
812 117
812 183
1 0 29 0 0 4096 0 9 0 0 139 2
792 117
792 192
1 0 28 0 0 4096 0 10 0 0 138 2
772 117
772 201
1 0 27 0 0 4096 0 11 0 0 137 2
752 117
752 210
2 0 29 0 0 0 0 17 0 0 139 2
718 123
718 192
3 0 28 0 0 0 0 17 0 0 138 2
712 123
712 201
4 0 27 0 0 0 0 17 0 0 137 4
706 123
706 205
707 205
707 210
1 0 34 0 0 0 0 13 0 0 144 2
656 118
656 136
1 0 33 0 0 0 0 14 0 0 143 2
636 118
636 145
1 0 32 0 0 0 0 15 0 0 142 2
616 118
616 154
1 0 31 0 0 0 0 16 0 0 141 2
596 118
596 163
1 0 34 0 0 0 0 18 0 0 144 2
570 122
570 136
2 0 33 0 0 0 0 18 0 0 143 2
564 122
564 145
3 0 32 0 0 0 0 18 0 0 142 2
558 122
558 154
4 0 31 0 0 0 0 18 0 0 141 2
552 122
552 163
0 0 35 0 0 12672 0 0 0 0 0 5
821 130
821 170
858 170
858 126
820 126
0 0 10 0 0 4480 0 0 0 0 0 2
59 640
773 640
0 0 9 0 0 4480 0 0 0 0 0 2
59 656
772 656
0 0 36 0 0 8576 0 0 0 0 0 5
658 488
696 488
696 532
658 532
658 488
0 0 37 0 0 12672 0 0 0 0 0 5
659 438
659 481
696 481
696 434
658 434
0 0 38 0 0 8576 0 0 0 0 0 5
659 382
696 382
696 426
659 426
659 382
0 0 39 0 0 4480 0 0 0 0 0 5
659 322
659 373
695 373
695 322
659 322
0 0 14 0 0 4224 0 0 0 0 0 2
84 365
669 365
0 0 24 0 0 4224 0 0 0 0 0 2
85 355
670 355
0 0 25 0 0 4224 0 0 0 0 0 2
84 345
669 345
0 0 26 0 0 4224 0 0 0 0 0 2
83 335
668 335
0 0 11 0 0 4224 0 0 0 0 0 2
85 473
670 473
0 0 20 0 0 4224 0 0 0 0 0 2
86 463
671 463
0 0 19 0 0 4224 0 0 0 0 0 2
85 453
670 453
0 0 18 0 0 4224 0 0 0 0 0 2
84 443
669 443
0 0 12 0 0 4224 0 0 0 0 0 2
87 524
672 524
0 0 17 0 0 4224 0 0 0 0 0 2
88 514
673 514
0 0 16 0 0 4224 0 0 0 0 0 2
87 504
672 504
0 0 15 0 0 4224 0 0 0 0 0 2
86 494
671 494
0 0 13 0 0 4224 0 0 0 0 0 2
87 419
672 419
0 0 23 0 0 4224 0 0 0 0 0 2
88 409
673 409
0 0 22 0 0 4224 0 0 0 0 0 2
87 399
672 399
0 0 21 0 0 4224 0 0 0 0 0 2
86 389
671 389
0 0 8 0 0 4224 0 0 0 0 0 2
14 716
987 716
0 0 7 0 0 4224 0 0 0 0 0 2
14 705
988 705
0 0 6 0 0 4224 0 0 0 0 0 2
14 694
987 694
0 0 5 0 0 4224 0 0 0 0 0 2
14 684
988 684
0 0 27 0 0 4224 0 0 0 0 0 2
15 210
836 210
0 0 28 0 0 4224 0 0 0 0 0 2
14 201
836 201
0 0 29 0 0 4224 0 0 0 0 0 2
15 192
836 192
0 0 30 0 0 4224 0 0 0 0 0 2
15 183
837 183
0 0 31 0 0 4224 0 0 0 0 0 2
13 163
834 163
0 0 32 0 0 4224 0 0 0 0 0 2
12 154
834 154
0 0 33 0 0 4224 0 0 0 0 0 2
13 145
834 145
0 0 34 0 0 4224 0 0 0 0 0 2
13 136
835 136
18
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
696 320 737 344
700 324 732 340
4 BusW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
698 380 739 404
702 384 734 400
4 BusX
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
698 431 739 455
702 435 734 451
4 BusY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
698 484 739 508
702 488 734 504
4 BusZ
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
698 340 731 364
702 344 726 360
3 Add
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
695 400 752 424
699 404 747 420
6 Buffer
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
698 451 739 475
702 455 734 471
4 Nand
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
698 501 731 525
702 505 726 521
3 Sub
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1017 694 1058 718
1021 698 1053 714
4 BusU
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
858 140 899 164
862 144 894 160
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
859 190 900 214
863 194 895 210
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
663 31 704 55
667 35 699 51
4 In`s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 7
707 543 772 567
711 547 767 563
7 Funcoes
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
890 569 939 593
894 573 934 589
5 Out`s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 20
756 326 797 430
760 330 792 410
20 Dec.
 0
 1
 2
 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 98
799 327 1000 431
803 331 995 411
98 S1  S0    BusU
 0   0    BusA+BusB
 0   1    BusA
 1   0    BusA.BusB(neg)
 1   1    BusA-BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
811 284 852 328
815 288 847 320
10 Ctrl
In`s
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 14
900 283 965 327
904 287 960 319
14 Funcoes
Out`s
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
