CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
8912914 0
0
6 Title:
5 Name:
0
0
0
14
9 2-In AND~
219 285 345 0 1 22
0 0
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 2 0
1 U
3976 0 0
2
45193.1 0
0
9 2-In AND~
219 285 309 0 1 22
0 0
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 2 0
1 U
7634 0 0
2
45193.1 0
0
9 2-In AND~
219 285 274 0 1 22
0 0
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
523 0 0
2
45193.1 0
0
9 2-In AND~
219 286 239 0 1 22
0 0
0
0 0 96 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
6748 0 0
2
45193.1 0
0
9 Inverter~
13 232 190 0 1 22
0 0
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1B
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
6901 0 0
2
45193.1 0
0
9 Inverter~
13 208 189 0 1 22
0 0
0
0 0 96 270
6 74LS04
-21 -19 21 -11
3 U1A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
842 0 0
2
45193.1 0
0
14 Logic Display~
6 602 133 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 M1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3277 0 0
2
45193.1 3
0
14 Logic Display~
6 582 133 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 M2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4212 0 0
2
45193.1 2
0
14 Logic Display~
6 562 133 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 M3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4720 0 0
2
45193.1 1
0
14 Logic Display~
6 622 133 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 M0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5551 0 0
2
45193.1 0
0
14 Logic Display~
6 184 132 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 S0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6986 0 0
2
45193.1 1
0
14 Logic Display~
6 164 132 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 S1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8745 0 0
2
45193.1 0
0
8 Hex Key~
166 131 127 0 11 12
0 0 0 0 0 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
9592 0 0
2
45193.1 0
0
12 Hex Display~
7 657 128 0 16 19
10 0 0 0 0 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
8748 0 0
2
45193.1 0
0
36
0 0 0 0 0 32 0 0 0 0 0 2
672 84
552 84
0 0 0 0 0 32 0 0 0 0 0 2
114 83
192 83
0 0 0 0 0 32 0 0 0 0 0 2
659 254
872 254
0 0 0 0 0 32 0 0 0 0 0 2
699 234
699 324
0 0 0 0 0 32 0 0 0 0 0 2
758 234
758 324
0 0 0 0 0 32 0 0 0 0 0 5
659 234
872 234
872 324
659 324
659 234
0 0 0 0 0 256 0 0 0 0 0 5
152 149
635 149
635 404
152 404
152 149
3 0 0 0 0 0 0 1 0 0 34 2
306 345
562 345
3 0 0 0 0 0 0 2 0 0 33 2
306 309
582 309
3 0 0 0 0 0 0 3 0 0 32 2
306 274
602 274
3 0 0 0 0 0 0 4 0 0 31 2
307 239
622 239
2 0 0 0 0 0 0 1 0 0 35 2
261 354
184 354
1 0 0 0 0 0 0 1 0 0 36 2
261 336
164 336
2 0 0 0 0 256 0 2 0 0 21 2
261 318
235 318
1 0 0 0 0 0 0 2 0 0 36 2
261 300
164 300
2 0 0 0 0 0 0 3 0 0 35 2
261 283
184 283
1 0 0 0 0 256 0 3 0 0 20 2
261 265
211 265
2 0 0 0 0 256 0 4 0 0 21 2
262 248
235 248
1 0 0 0 0 256 0 4 0 0 20 2
262 230
211 230
2 0 0 0 0 256 0 6 0 0 0 2
211 207
211 389
2 0 0 0 0 256 0 5 0 0 0 2
235 208
235 389
4 0 0 0 0 0 0 14 0 0 34 3
648 152
648 169
562 169
3 0 0 0 0 0 0 14 0 0 33 3
654 152
654 180
582 180
2 0 0 0 0 0 0 14 0 0 32 3
660 152
660 191
602 191
1 0 0 0 0 0 0 14 0 0 31 3
666 152
666 201
622 201
2 0 0 0 0 0 0 13 0 0 36 3
134 151
134 200
164 200
1 0 0 0 0 0 0 13 0 0 35 3
140 151
140 188
184 188
0 1 0 0 0 0 0 0 5 35 0 3
184 156
235 156
235 172
0 1 0 0 0 0 0 0 6 36 0 3
164 166
211 166
211 171
1 0 0 0 0 0 0 5 0 0 0 3
235 172
235 170
246 170
1 0 0 0 0 0 0 10 0 0 0 2
622 151
622 391
1 0 0 0 0 0 0 7 0 0 0 2
602 151
602 391
1 0 0 0 0 0 0 8 0 0 0 2
582 151
582 391
1 0 0 0 0 0 0 9 0 0 0 2
562 151
562 391
1 0 0 0 0 0 0 11 0 0 0 2
184 150
184 391
1 0 0 0 0 0 0 12 0 0 0 2
164 150
164 391
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
586 61 639 85
592 65 632 81
5 Out's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
130 60 175 84
136 64 168 80
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
339 124 432 148
345 128 425 144
10 Decode2bit
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 105
699 235 872 339
705 239 865 319
105 S1 S0    M3 M2 M1 M0
0  0     0  0  0  1
0  1     0  0  1  0 
1  0     0  1  0  0
1  1     1  0  0  0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
658 233 703 337
664 237 696 317
16 Dec.
0
1
2
3
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
