CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
13
12 Hex Display~
7 779 196 0 18 19
10 3 2 11 12 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
5130 0 0
2
5.90094e-315 5.40342e-315
0
14 Logic Display~
6 337 188 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 A
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
391 0 0
2
5.90094e-315 5.39824e-315
0
14 Logic Display~
6 360 188 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 B
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
5.90094e-315 5.39306e-315
0
14 Logic Display~
6 383 188 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Te
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.90094e-315 5.38788e-315
0
14 Logic Display~
6 724 183 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
1 W
-4 -21 3 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.90094e-315 5.37752e-315
0
14 Logic Display~
6 699 183 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Ts
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.90094e-315 5.36716e-315
0
9 2-In XOR~
219 507 265 0 3 22
0 4 9 3
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
8901 0 0
2
5.90094e-315 5.3568e-315
0
9 2-In XOR~
219 421 325 0 3 22
0 6 5 9
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
7361 0 0
2
5.90094e-315 5.34643e-315
0
9 2-In AND~
219 517 391 0 3 22
0 9 4 7
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4747 0 0
2
5.90094e-315 5.32571e-315
0
8 2-In OR~
219 610 466 0 3 22
0 7 8 2
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U2A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
972 0 0
2
5.90094e-315 5.30499e-315
0
9 2-In AND~
219 434 470 0 3 22
0 6 5 8
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3472 0 0
2
5.90094e-315 5.26354e-315
0
8 Hex Key~
166 279 184 0 11 12
0 13 14 15 16 0 0 0 0 0
4 52
0
0 0 4640 0
0
4 KPD1
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9998 0 0
2
5.90094e-315 0
0
10 MT.Add1bit
94 524 519 0 1 11
0 0
10 MT.Add1bit
1 0 4736 0
0
2 U4
68 -36 82 -28
0
0
0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 0 0 0 0
1 U
3536 0 0
2
45193.8 0
0
35
2 0 2 0 0 12288 0 13 0 0 32 7
460 520
460 521
456 521
456 565
694 565
694 516
699 516
1 0 3 0 0 8192 0 13 0 0 31 5
524 544
524 554
719 554
719 525
724 525
3 0 4 0 0 12288 0 13 0 0 33 7
594 519
594 520
598 520
598 550
388 550
388 524
383 524
5 0 5 0 0 8192 0 13 0 0 34 5
559 486
559 483
449 483
449 512
360 512
4 0 6 0 0 16384 0 13 0 0 35 5
496 486
496 477
459 477
459 500
337 500
0 0 1 0 0 4128 0 0 0 0 0 2
824 288
1068 288
0 0 1 0 0 32 0 0 0 0 0 5
820 465
1030 465
1030 506
820 506
820 465
0 0 1 0 0 32 0 0 0 0 0 2
1018 264
1018 423
0 0 1 0 0 32 0 0 0 0 0 2
948 264
948 423
0 0 1 0 0 32 0 0 0 0 0 2
869 264
869 423
0 0 1 0 0 32 0 0 0 0 0 5
824 264
1068 264
1068 423
824 423
824 264
0 0 1 0 0 4256 0 0 0 0 0 2
327 360
736 360
2 0 2 0 0 0 0 1 0 0 32 3
782 220
782 238
699 238
1 0 3 0 0 0 0 1 0 0 31 3
788 220
788 248
724 248
0 0 6 0 0 0 0 0 0 0 35 3
276 225
276 246
337 246
0 0 5 0 0 0 0 0 0 0 34 3
282 225
282 234
360 234
0 0 4 0 0 0 0 0 0 0 33 2
288 225
383 225
3 0 2 0 0 0 0 10 0 0 32 2
643 466
699 466
3 0 3 0 0 0 0 7 0 0 31 2
540 265
724 265
3 1 7 0 0 8320 0 9 10 0 0 4
538 391
590 391
590 457
597 457
3 2 8 0 0 4224 0 11 10 0 0 4
455 470
588 470
588 475
597 475
2 0 5 0 0 0 0 11 0 0 34 2
410 479
360 479
1 0 6 0 0 0 0 11 0 0 35 2
410 461
337 461
2 0 4 0 0 0 0 9 0 0 33 2
493 400
383 400
2 0 5 0 0 0 0 8 0 0 34 2
405 334
360 334
1 0 6 0 0 0 0 8 0 0 35 2
405 316
337 316
0 1 9 0 0 4480 0 0 9 28 0 3
480 325
480 382
493 382
3 2 9 0 0 0 0 8 7 0 0 4
454 325
481 325
481 274
491 274
1 0 4 0 0 0 0 7 0 0 33 2
491 256
383 256
0 0 10 0 0 12672 0 0 0 0 0 5
321 204
746 204
746 561
316 561
316 204
1 0 3 0 0 4224 0 5 0 0 0 2
724 201
724 542
1 0 2 0 0 4224 0 6 0 0 0 2
699 201
699 543
1 0 4 0 0 4224 0 4 0 0 0 2
383 206
383 543
1 0 5 0 0 4224 0 3 0 0 0 2
360 206
360 544
1 0 6 0 0 4224 0 2 0 0 0 2
337 206
337 545
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 63
875 268 936 452
881 272 929 416
63 A B Te
0 0 0 
0 0 1
0 1 0
0 1 1
1 0 0
1 0 1
1 1 0
1 1 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 52
963 270 1008 454
969 274 1001 418
52 Ts W
0  0
0  1
0  1
1  0
0  1
1  0
1  0
1  1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
823 268 868 292
829 271 861 287
4 Dec.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1023 268 1068 292
1029 272 1061 288
4 Dec.
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
835 286 856 450
841 290 849 418
22 0
1
2
3
4
5
6
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 22
1033 288 1054 452
1039 292 1047 420
22 0
1
2
3
4
5
6
7
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 45
820 466 1033 510
826 470 1026 502
45 W = A (+) B (+) Te
Ts = A.B + Te . (A (+) B)
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
