CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
8912914 0
0
6 Title:
5 Name:
0
0
0
14
14 Logic Display~
6 738 281 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3835 0 0
2
45192.7 3
0
14 Logic Display~
6 757 281 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3670 0 0
2
45192.7 2
0
14 Logic Display~
6 777 281 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5616 0 0
2
45192.7 1
0
14 Logic Display~
6 797 281 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 X0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9323 0 0
2
45192.7 0
0
7 Buffer~
58 511 268 0 1 22
0 0
0
0 0 608 270
4 4050
-14 -19 14 -11
3 U1D
13 -5 34 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 4 1 0
1 U
317 0 0
2
45192.7 0
0
7 Buffer~
58 458 268 0 1 22
0 0
0
0 0 608 270
4 4050
-14 -19 14 -11
3 U1C
13 -5 34 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 3 1 0
1 U
3108 0 0
2
45192.7 0
0
7 Buffer~
58 407 268 0 1 22
0 0
0
0 0 608 270
4 4050
-14 -19 14 -11
3 U1B
13 -5 34 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 2 1 0
1 U
4299 0 0
2
45192.7 0
0
7 Buffer~
58 354 267 0 1 22
0 0
0
0 0 608 270
4 4050
-14 -19 14 -11
3 U1A
13 -5 34 3
0
14 DVCC=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 0 0
65 0 0 0 6 1 1 0
1 U
9672 0 0
2
45192.7 0
0
14 Logic Display~
6 208 136 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7876 0 0
2
45192.7 0
0
14 Logic Display~
6 188 136 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6369 0 0
2
45192.7 0
0
14 Logic Display~
6 168 136 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9172 0 0
2
45192.7 0
0
14 Logic Display~
6 149 136 0 1 2
10 0
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7100 0 0
2
45192.7 0
0
12 Hex Display~
7 834 284 0 16 19
10 0 0 0 0 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusX
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3820 0 0
2
45192.7 0
0
8 Hex Key~
166 116 133 0 11 12
0 0 0 0 0 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 0 0 0 0 0
3 KPD
7678 0 0
2
45192.7 0
0
37
0 0 0 0 0 32 0 0 0 0 0 2
851 239
729 239
0 0 0 0 0 32 0 0 0 0 0 2
98 92
216 92
1 0 0 0 0 0 0 13 0 0 33 2
843 308
843 319
2 0 0 0 0 0 0 13 0 0 32 2
837 308
837 330
3 0 0 0 0 0 0 13 0 0 31 2
831 308
831 340
4 0 0 0 0 0 0 13 0 0 30 2
825 308
825 351
1 0 0 0 0 0 0 1 0 0 30 2
738 299
738 351
1 0 0 0 0 0 0 2 0 0 31 2
757 299
757 340
1 0 0 0 0 0 0 3 0 0 32 2
777 299
777 330
1 0 0 0 0 0 0 4 0 0 33 2
797 299
797 319
0 0 0 0 0 256 0 0 0 0 0 5
330 167
330 369
561 369
561 163
330 163
0 0 0 0 0 272 0 0 0 0 0 5
908 310
942 310
942 364
908 364
908 310
0 0 0 0 0 256 0 0 0 0 0 5
25 173
59 173
59 227
25 227
25 173
2 0 0 0 0 0 0 5 0 0 33 2
511 283
511 319
1 0 0 0 0 0 0 5 0 0 37 2
511 253
511 182
2 0 0 0 0 0 0 6 0 0 32 2
458 283
458 330
1 0 0 0 0 0 0 6 0 0 36 2
458 253
458 193
2 0 0 0 0 0 0 7 0 0 31 2
407 283
407 340
1 0 0 0 0 0 0 7 0 0 35 2
407 253
407 204
2 0 0 0 0 0 0 8 0 0 30 2
354 282
354 351
1 0 0 0 0 0 0 8 0 0 34 2
354 252
354 215
1 0 0 0 0 0 0 9 0 0 37 2
208 154
208 182
1 0 0 0 0 0 0 10 0 0 36 2
188 154
188 193
1 0 0 0 0 0 0 11 0 0 35 2
168 154
168 204
1 0 0 0 0 0 0 12 0 0 34 2
149 154
149 215
1 0 0 0 0 0 0 14 0 0 37 2
125 157
125 182
2 0 0 0 0 0 0 14 0 0 36 2
119 157
119 193
3 0 0 0 0 0 0 14 0 0 35 2
113 157
113 204
4 0 0 0 0 0 0 14 0 0 34 2
107 157
107 215
0 0 0 0 0 0 0 0 0 0 0 2
43 351
929 351
0 0 0 0 0 0 0 0 0 0 0 2
43 340
929 340
0 0 0 0 0 0 0 0 0 0 0 2
42 330
928 330
0 0 0 0 0 0 0 0 0 0 0 2
42 319
928 319
0 0 0 0 0 0 0 0 0 0 0 2
41 215
576 215
0 0 0 0 0 0 0 0 0 0 0 2
40 204
576 204
0 0 0 0 0 0 0 0 0 0 0 2
39 193
576 193
0 0 0 0 0 0 0 0 0 0 0 2
39 182
576 182
5
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
764 215 817 239
770 219 810 235
5 Out's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
134 67 179 111
140 71 172 103
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
901 289 946 313
907 293 939 309
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
19 152 64 176
25 156 57 172
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
404 139 505 163
410 143 498 159
11 Buffer.4bit
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
