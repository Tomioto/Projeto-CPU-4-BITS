CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
100 C:\Users\Matheus Mioto\OneDrive - UNIRP\Desktop\Arquivos faculdade\CircuitMaker\CircuitMaker\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9961490 0
0
6 Title:
5 Name:
0
0
0
20
12 Hex Display~
7 1043 447 0 16 19
10 6 7 8 9 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 BusY
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5130 0 0
2
5.90094e-315 5.43451e-315
0
14 Logic Display~
6 200 74 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
391 0 0
2
5.90094e-315 5.43192e-315
0
14 Logic Display~
6 222 74 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3124 0 0
2
5.90094e-315 5.42933e-315
0
14 Logic Display~
6 245 74 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3421 0 0
2
5.90094e-315 5.42414e-315
0
14 Logic Display~
6 266 74 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 A0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8157 0 0
2
5.90094e-315 5.41896e-315
0
14 Logic Display~
6 386 72 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.90094e-315 5.41378e-315
0
14 Logic Display~
6 406 72 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.90094e-315 5.4086e-315
0
14 Logic Display~
6 427 72 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.90094e-315 5.40342e-315
0
14 Logic Display~
6 448 72 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 B0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.90094e-315 5.39824e-315
0
14 Logic Display~
6 985 432 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y0
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.90094e-315 5.39306e-315
0
14 Logic Display~
6 964 432 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.90094e-315 5.38788e-315
0
14 Logic Display~
6 943 432 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.90094e-315 5.37752e-315
0
14 Logic Display~
6 923 432 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 Y3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.90094e-315 5.36716e-315
0
10 2-In NAND~
219 599 398 0 3 22
0 2 10 9
0
0 0 96 270
6 74LS00
-14 -24 28 -16
3 U1D
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
4597 0 0
2
5.90094e-315 5.3568e-315
0
10 2-In NAND~
219 642 397 0 3 22
0 3 11 8
0
0 0 96 270
6 74LS00
-14 -24 28 -16
3 U1C
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3835 0 0
2
5.90094e-315 5.34643e-315
0
10 2-In NAND~
219 683 397 0 3 22
0 4 12 7
0
0 0 96 270
6 74LS00
-14 -24 28 -16
3 U1B
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3670 0 0
2
5.90094e-315 5.32571e-315
0
10 2-In NAND~
219 724 397 0 3 22
0 5 13 6
0
0 0 96 270
6 74LS00
-14 -24 28 -16
3 U1A
19 -7 40 1
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
5616 0 0
2
5.90094e-315 5.30499e-315
0
8 Hex Key~
166 326 82 0 11 12
0 19 20 21 22 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusB
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
9323 0 0
2
5.90094e-315 5.26354e-315
0
8 Hex Key~
166 159 81 0 11 12
0 23 24 25 26 0 0 0 0 0
0 48
0
0 0 4640 0
0
4 BusA
-14 -34 14 -26
0
0
0
0
0
4 SIP4
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
3 KPD
317 0 0
2
5.90094e-315 0
0
12 MT.Nand4bits
94 295 390 0 1 25
0 0
12 MT.Nand4bits
1 0 4736 0
0
2 U2
42 1 56 9
0
0
0
0
0
0
25

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0 0 0 0 0
1 U
3108 0 0
2
45193.9 0
0
70
9 0 2 0 0 4096 0 20 0 0 67 2
295 366
295 308
10 0 3 0 0 4096 0 20 0 0 68 2
304 366
304 295
11 0 4 0 0 4096 0 20 0 0 69 2
313 366
313 281
12 0 5 0 0 4096 0 20 0 0 70 2
322 366
322 267
4 0 6 0 0 4096 0 20 0 0 46 4
322 425
322 480
356 480
356 495
3 0 7 0 0 4096 0 20 0 0 44 4
304 425
304 492
338 492
338 507
2 0 8 0 0 4096 0 20 0 0 45 4
268 425
268 505
302 505
302 520
1 0 9 0 0 4096 0 20 0 0 43 4
251 425
251 518
285 518
285 533
5 0 10 0 0 4096 0 20 0 0 63 2
250 366
250 202
6 0 11 0 0 4096 0 20 0 0 64 2
260 366
260 189
7 0 12 0 0 4096 0 20 0 0 65 2
269 366
269 175
8 0 13 0 0 4096 0 20 0 0 66 2
278 366
278 161
0 0 14 0 0 4224 0 0 0 0 0 2
690 76
779 76
3 0 6 0 0 4096 0 17 0 0 46 2
725 423
725 495
3 0 7 0 0 4096 0 16 0 0 44 2
684 423
684 507
3 0 8 0 0 4096 0 15 0 0 45 2
643 423
643 520
3 0 9 0 0 4096 0 14 0 0 43 2
600 424
600 533
0 0 15 0 0 12672 0 0 0 0 0 6
26 257
26 321
82 321
82 251
26 251
26 257
0 0 16 0 0 12672 0 0 0 0 0 6
26 153
26 217
82 217
82 147
26 147
26 153
0 0 1 0 0 4128 0 0 0 0 0 2
624 43
624 104
0 0 1 0 0 4128 0 0 0 0 0 2
522 66
794 66
0 0 1 0 0 32 0 0 0 0 0 5
522 43
794 43
794 104
522 104
522 43
0 0 17 0 0 12672 0 0 0 0 0 5
500 142
500 553
777 553
777 138
500 138
1 0 5 0 0 4096 0 17 0 0 70 2
734 372
734 267
2 0 13 0 0 4096 0 17 0 0 66 2
716 372
716 161
1 0 4 0 0 0 0 16 0 0 69 4
693 372
693 296
670 296
670 281
2 0 12 0 0 0 0 16 0 0 65 4
675 372
675 190
652 190
652 175
1 0 3 0 0 0 0 15 0 0 68 4
652 372
652 310
607 310
607 295
2 0 11 0 0 0 0 15 0 0 64 4
634 372
634 204
589 204
589 189
1 0 2 0 0 8192 0 14 0 0 67 4
609 373
609 323
540 323
540 308
2 0 10 0 0 0 0 14 0 0 63 4
591 373
591 217
522 217
522 202
0 0 1 0 0 32 0 0 0 0 0 2
912 401
1061 401
0 0 1 0 0 4256 0 0 0 0 0 2
142 45
458 45
1 0 6 0 0 0 0 1 0 0 46 2
1052 471
1052 495
2 0 7 0 0 0 0 1 0 0 44 2
1046 471
1046 507
3 0 8 0 0 0 0 1 0 0 45 2
1040 471
1040 520
4 0 9 0 0 0 0 1 0 0 43 2
1034 471
1034 533
1 0 6 0 0 0 0 10 0 0 46 2
985 450
985 495
1 0 7 0 0 0 0 11 0 0 44 2
964 450
964 507
1 0 8 0 0 0 0 12 0 0 45 2
943 450
943 520
1 0 9 0 0 0 0 13 0 0 43 2
923 450
923 533
0 0 18 0 0 12672 0 0 0 0 0 6
1080 484
1080 548
1137 548
1137 475
1080 475
1080 484
0 0 9 0 0 4224 0 0 0 0 0 2
55 533
1111 533
0 0 7 0 0 4224 0 0 0 0 0 2
56 507
1112 507
0 0 8 0 0 4224 0 0 0 0 0 2
57 520
1111 520
0 0 6 0 0 4224 0 0 0 0 0 2
56 495
1112 495
1 0 5 0 0 4096 0 9 0 0 70 2
448 90
448 267
1 0 4 0 0 4096 0 8 0 0 69 2
427 90
427 281
1 0 3 0 0 4096 0 7 0 0 68 2
406 90
406 295
1 0 2 0 0 4096 0 6 0 0 67 2
386 90
386 308
0 0 13 0 0 0 0 0 0 0 66 2
336 110
336 161
0 0 12 0 0 0 0 0 0 0 65 2
330 110
330 175
0 0 11 0 0 0 0 0 0 0 64 2
324 110
324 189
0 0 10 0 0 0 0 0 0 0 63 2
318 110
318 202
1 0 13 0 0 0 0 5 0 0 66 2
266 92
266 161
1 0 12 0 0 0 0 4 0 0 65 2
245 92
245 175
1 0 11 0 0 0 0 3 0 0 64 2
222 92
222 189
1 0 10 0 0 0 0 2 0 0 63 2
200 92
200 202
0 0 13 0 0 0 0 0 0 0 66 2
168 110
168 161
0 0 12 0 0 0 0 0 0 0 65 2
162 110
162 175
0 0 11 0 0 0 0 0 0 0 64 2
156 110
156 189
0 0 10 0 0 0 0 0 0 0 63 2
150 110
150 202
0 0 10 0 0 4224 0 0 0 0 0 2
53 202
936 202
0 0 11 0 0 4224 0 0 0 0 0 2
54 189
936 189
0 0 12 0 0 4224 0 0 0 0 0 2
54 175
937 175
0 0 13 0 0 4224 0 0 0 0 0 2
52 161
938 161
0 0 2 0 0 4224 0 0 0 0 0 2
54 308
937 308
0 0 3 0 0 4224 0 0 0 0 0 2
55 295
937 295
0 0 4 0 0 4224 0 0 0 0 0 2
55 281
938 281
0 0 5 0 0 4224 0 0 0 0 0 2
53 267
939 267
8
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
591 20 684 44
597 24 677 40
10 Nand.4bits
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
590 114 683 138
596 118 676 134
10 Nand.4bits
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 60
520 44 789 108
526 48 782 96
60    In's            Out's

 BusA, BusB   BusY = BusA . BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
1079 452 1124 476
1085 456 1117 472
4 BusY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
31 123 76 147
37 127 69 143
4 BusA
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
33 229 78 253
39 233 71 249
4 BusB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 4
265 21 310 45
271 25 303 41
4 In's
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
959 377 1012 401
965 381 1005 397
5 Out's
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
